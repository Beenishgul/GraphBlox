`define IOB_CACHE_LRU 0
`define IOB_CACHE_PLRU_MRU 1
`define IOB_CACHE_PLRU_TREE 2
`define IOB_CACHE_WRITE_THROUGH 0
`define IOB_CACHE_WRITE_BACK 1
`define IOB_CACHE_ADDR_W `IOB_CACHE_SWREG_ADDR_W
`define IOB_CACHE_DATA_W 32
`define IOB_CACHE_FE_ADDR_W 24
`define IOB_CACHE_FE_DATA_W 32
`define IOB_CACHE_BE_ADDR_W 24
`define IOB_CACHE_BE_DATA_W 512
`define IOB_CACHE_NWAYS_W 1
`define IOB_CACHE_NLINES_W 7
`define IOB_CACHE_WORD_OFFSET_W 3
`define IOB_CACHE_WTBUF_DEPTH_W 4
`define IOB_CACHE_REP_POLICY 0
`define IOB_CACHE_WRITE_POL 0 
`define IOB_CACHE_USE_CTRL 0
`define IOB_CACHE_USE_CTRL_CNT 0
`define IOB_CACHE_AXI NA
`define IOB_CACHE_AXI_ID_W 1
`define IOB_CACHE_AXI_LEN_W 4
`define IOB_CACHE_AXI_ID 0
`define IOB_CACHE_VERSION 16'h0010
