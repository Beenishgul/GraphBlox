    parameter ID_CU           = 0,
// --------------------------------------------------------------------------------------
// CU SETTINGS
// --------------------------------------------------------------------------------------
`include "topology_parameters.vh"
