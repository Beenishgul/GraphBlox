parameter NUM_CUS     = 1;
parameter NUM_BUNDLES = 4;
parameter NUM_LANES   = 4;
parameter NUM_ENGINES = 2;
parameter NUM_MODULES = 3;
parameter NUM_CHANNELS           = 2;
parameter CACHE_CONFIG_MAX_NUM_WAYS   = 4;
parameter CACHE_CONFIG_MAX_SIZE = 32768;

parameter NUM_CHANNELS_WIDTH_BITS = 2;
parameter NUM_CUS_WIDTH_BITS      = 1;
parameter NUM_BUNDLES_WIDTH_BITS  = 4;
parameter NUM_LANES_WIDTH_BITS    = 4;
parameter NUM_ENGINES_WIDTH_BITS  = 2;
parameter NUM_MODULES_WIDTH_BITS  = 3;
parameter CU_PACKET_SEQUENCE_ID_WIDTH_BITS = $clog2((96*NUM_BUNDLES)+(8*NUM_BUNDLES));
parameter BUFFER_0_WIDTH_BITS = 64;
parameter BUFFER_1_WIDTH_BITS = 64;
parameter BUFFER_2_WIDTH_BITS = 64;
parameter BUFFER_3_WIDTH_BITS = 64;
parameter BUFFER_4_WIDTH_BITS = 64;
parameter BUFFER_5_WIDTH_BITS = 64;
parameter BUFFER_6_WIDTH_BITS = 64;
parameter BUFFER_7_WIDTH_BITS = 64;
parameter BUFFER_8_WIDTH_BITS = 64;
parameter BUFFER_9_WIDTH_BITS = 64;
