.CU_BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY (CU_BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY          ),
.CU_BUNDLES_CONFIG_MAX_CAST_WIDTH_ARRAY  (CU_BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY          ),
.CU_BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY  (CU_BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY ),
.CU_BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY (CU_BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY),
.CU_BUNDLES_CONFIG_ARRAY                 (CU_BUNDLES_CONFIG_ARRAY                          ),
.CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN  (CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN           ),       
.CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH(CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH         ),  
.CU_BUNDLES_CONFIG_CAST_WIDTH_ARRAY      (CU_BUNDLES_CONFIG_CAST_WIDTH_ARRAY               ),
.CU_BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY (CU_BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY          ),
.CU_BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY(CU_BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY         ),
.CU_BUNDLES_CONFIG_MERGE_CONNECT_ARRAY   (CU_BUNDLES_CONFIG_MERGE_CONNECT_ARRAY            ),
.CU_BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY(CU_BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY ),
.CU_BUNDLES_CONFIG_MERGE_WIDTH_ARRAY     (CU_BUNDLES_CONFIG_MERGE_WIDTH_ARRAY              ),
.CU_BUNDLES_COUNT_ARRAY                  (CU_BUNDLES_COUNT_ARRAY                           ),
.CU_BUNDLES_ENGINE_ID_ARRAY              (CU_BUNDLES_ENGINE_ID_ARRAY                       ),
.CU_BUNDLES_LANES_COUNT_ARRAY            (CU_BUNDLES_LANES_COUNT_ARRAY                     ),
.CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY    (CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY             ),
.BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY    (BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY             ),
.BUNDLES_CONFIG_MAX_CAST_WIDTH_ARRAY     (BUNDLES_CONFIG_MAX_CAST_WIDTH_ARRAY              ),
.BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY    (BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY     ),
.BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY   (BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY    ),
.BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY   (BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY    ),
.BUNDLES_CONFIG_ARRAY                    (BUNDLES_CONFIG_ARRAY                             ),
.BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN     (BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN              ),        
.BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH   (BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH            ),  
.BUNDLES_CONFIG_CAST_WIDTH_ARRAY         (BUNDLES_CONFIG_CAST_WIDTH_ARRAY                  ),
.BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY    (BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY             ),
.BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY   (BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY            ),
.BUNDLES_CONFIG_MERGE_CONNECT_ARRAY      (BUNDLES_CONFIG_MERGE_CONNECT_ARRAY               ),
.BUNDLES_CONFIG_MERGE_WIDTH_ARRAY        (BUNDLES_CONFIG_MERGE_WIDTH_ARRAY                 ),
.BUNDLES_ENGINE_ID_ARRAY                 (BUNDLES_ENGINE_ID_ARRAY                          ),
.LANES_CONFIG_MAX_MERGE_WIDTH_ARRAY      (LANES_CONFIG_MAX_MERGE_WIDTH_ARRAY               ),
.LANES_CONFIG_MAX_CAST_WIDTH_ARRAY       (LANES_CONFIG_MAX_CAST_WIDTH_ARRAY                ),
.LANES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY  (LANES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY           ),
.LANES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY (LANES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY          ),
.LANES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY (LANES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY          ),
.LANES_CONFIG_ARRAY                      (LANES_CONFIG_ARRAY                               ),
.LANES_CONFIG_ARRAY_ENGINE_SEQ_MIN       (LANES_CONFIG_ARRAY_ENGINE_SEQ_MIN                ),             
.LANES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH     (LANES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH              ),
.LANES_CONFIG_CAST_WIDTH_ARRAY           (LANES_CONFIG_CAST_WIDTH_ARRAY                    ),
.LANES_CONFIG_LANE_CAST_WIDTH_ARRAY      (LANES_CONFIG_LANE_CAST_WIDTH_ARRAY               ),
.LANES_CONFIG_LANE_MERGE_WIDTH_ARRAY     (LANES_CONFIG_LANE_MERGE_WIDTH_ARRAY              ),
.LANES_CONFIG_MERGE_CONNECT_ARRAY        (LANES_CONFIG_MERGE_CONNECT_ARRAY                 ),
.LANES_CONFIG_MERGE_WIDTH_ARRAY          (LANES_CONFIG_MERGE_WIDTH_ARRAY                   ),
.LANES_COUNT_ARRAY                       (LANES_COUNT_ARRAY                                ),
.LANES_ENGINE_ID_ARRAY                   (LANES_ENGINE_ID_ARRAY                            ),
.LANES_ENGINES_COUNT_ARRAY               (LANES_ENGINES_COUNT_ARRAY                        ),
.ENGINES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY   (ENGINES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY    ),
.ENGINES_CONFIG_MAX_MERGE_WIDTH_ARRAY    (ENGINES_CONFIG_MAX_MERGE_WIDTH_ARRAY             ),
.ENGINES_CONFIG_MAX_CAST_WIDTH_ARRAY     (ENGINES_CONFIG_MAX_CAST_WIDTH_ARRAY              ),
.ENGINES_CONFIG                          (ENGINES_CONFIG_ARRAY[j]                          ),
.ENGINES_CONFIG_ARRAY                    (ENGINES_CONFIG_ARRAY                             ),
.ENGINES_CONFIG_ARRAY_ENGINE_SEQ_MIN     (ENGINES_CONFIG_ARRAY_ENGINE_SEQ_MIN              ),                      
.ENGINES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH   (ENGINES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH            ),  
.ENGINES_CONFIG_CAST_WIDTH_ARRAY         (ENGINES_CONFIG_CAST_WIDTH_ARRAY                  ),
.ENGINES_CONFIG_LANE_CAST_WIDTH_ARRAY    (ENGINES_CONFIG_LANE_CAST_WIDTH_ARRAY             ),
.ENGINES_CONFIG_LANE_MERGE_WIDTH_ARRAY   (ENGINES_CONFIG_LANE_MERGE_WIDTH_ARRAY            ),
.ENGINES_CONFIG_MERGE_CONNECT_ARRAY      (ENGINES_CONFIG_MERGE_CONNECT_ARRAY               ),
.ENGINES_CONFIG_MERGE_WIDTH_ARRAY        (ENGINES_CONFIG_MERGE_WIDTH_ARRAY                 ),
.ENGINES_COUNT_ARRAY                     (ENGINES_COUNT_ARRAY                              ),
.ENGINES_ENGINE_ID_ARRAY                 (ENGINES_ENGINE_ID_ARRAY                          ),
.ID_BUNDLE                               (ID_BUNDLE                                        ),
.ID_CU                                   (ID_CU                                            ),
.ID_ENGINE                               (j                                                ),
.ID_LANE                                 (ID_LANE                                          ),
.ID_RELATIVE                             (ENGINES_ENGINE_ID_ARRAY[j]                       ),
.LANE_CAST_WIDTH                         (LANE_CAST_WIDTH                                  ),
.LANE_MERGE_WIDTH                        (LANE_MERGE_WIDTH                                 ),
.ENGINE_CAST_WIDTH                       (ENGINES_CONFIG_CAST_WIDTH_ARRAY[j]               ),
.ENGINE_MERGE_WIDTH                      (ENGINES_CONFIG_MERGE_WIDTH_ARRAY[j]              ),
.NUM_BUNDLES                             (NUM_BUNDLES                                      ),
.NUM_ENGINES                             (NUM_ENGINES                                      ),
.FIFO_WRITE_DEPTH 					     (32                                               ),
.PROG_THRESH      						 (16                                               ),
.ENGINE_SEQ_WIDTH                        (ENGINES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH[j]         ),
.ENGINE_SEQ_MIN                          (ENGINES_CONFIG_ARRAY_ENGINE_SEQ_MIN[j]           ),
.NUM_LANES                               (NUM_LANES                                        )
