
    // Slave MM VIP instantiation
    import slv_m00_axi_vip_pkg::*;
        

    // Slave MM VIP instantiation
    import slv_m01_axi_vip_pkg::*;
        