// --------------------------------------------------------------------------------------
// CU SETTINGS
// --------------------------------------------------------------------------------------

`include "topology_parameters.vh"
