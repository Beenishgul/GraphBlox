
parameter integer C_M00_AXI_ADDR_WIDTH       = 64 ,
parameter integer C_M00_AXI_DATA_WIDTH       = 512 ,
parameter integer C_M00_AXI_ID_WIDTH         = 1   ,


parameter integer C_M01_AXI_ADDR_WIDTH       = 64 ,
parameter integer C_M01_AXI_DATA_WIDTH       = 512 ,
parameter integer C_M01_AXI_ID_WIDTH         = 1   ,

parameter integer C_S_AXI_CONTROL_ADDR_WIDTH = 12 ,
parameter integer C_S_AXI_CONTROL_DATA_WIDTH = 32