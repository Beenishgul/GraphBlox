
generate
     if(ID_BUNDLE == 0)
                    begin
                      assign lanes_fifo_request_cast_lane_out_signals_in[0][0]  = lanes_fifo_request_lane_out_signals_in[0];
                      assign lanes_fifo_request_lane_out_signals_out[0]         = lanes_fifo_request_cast_lane_out_signals_out [0][0];
                      assign lanes_fifo_response_lane_in_signals_out[0]         = lanes_fifo_response_merge_lane_in_signals_out[0][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][0] = lanes_fifo_response_lane_in_signals_in[0];
                      assign lanes_request_lane_out[0]                          = lanes_request_cast_lane_out[0][0];
                      assign lanes_response_merge_engine_in[0][0]               = lanes_response_engine_in[0];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][1].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][1]                                 = lanes_request_cast_lane_out[1][1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][1].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][2]                                 = lanes_request_cast_lane_out[2][1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][1].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][3].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][3].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][3]                                 = lanes_request_cast_lane_out[3][1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][0]  = lanes_fifo_request_lane_out_signals_in[1];
                      assign lanes_fifo_request_lane_out_signals_out[1]         = lanes_fifo_request_cast_lane_out_signals_out [1][0];
                      assign lanes_fifo_response_lane_in_signals_out[1]         = lanes_fifo_response_merge_lane_in_signals_out[1][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][0] = lanes_fifo_response_lane_in_signals_in[1];
                      assign lanes_request_lane_out[1]                          = lanes_request_cast_lane_out[1][0];
                      assign lanes_response_merge_engine_in[1][0]               = lanes_response_engine_in[1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][2].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][1]                                 = lanes_request_cast_lane_out[2][2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][2].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][2]                                 = lanes_request_cast_lane_out[3][2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][0]  = lanes_fifo_request_lane_out_signals_in[2];
                      assign lanes_fifo_request_lane_out_signals_out[2]         = lanes_fifo_request_cast_lane_out_signals_out [2][0];
                      assign lanes_fifo_response_lane_in_signals_out[2]         = lanes_fifo_response_merge_lane_in_signals_out[2][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][0] = lanes_fifo_response_lane_in_signals_in[2];
                      assign lanes_request_lane_out[2]                          = lanes_request_cast_lane_out[2][0];
                      assign lanes_response_merge_engine_in[2][0]               = lanes_response_engine_in[2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][3].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[2][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[2][1]                                 = lanes_request_cast_lane_out[3][3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][0]  = lanes_fifo_request_lane_out_signals_in[3];
                      assign lanes_fifo_request_lane_out_signals_out[3]         = lanes_fifo_request_cast_lane_out_signals_out [3][0];
                      assign lanes_fifo_response_lane_in_signals_out[3]         = lanes_fifo_response_merge_lane_in_signals_out[3][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[3][0] = lanes_fifo_response_lane_in_signals_in[3];
                      assign lanes_request_lane_out[3]                          = lanes_request_cast_lane_out[3][0];
                      assign lanes_response_merge_engine_in[3][0]               = lanes_response_engine_in[3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[4][0]  = lanes_fifo_request_lane_out_signals_in[4];
                      assign lanes_fifo_request_lane_out_signals_out[4]         = lanes_fifo_request_cast_lane_out_signals_out [4][0];
                      assign lanes_fifo_response_lane_in_signals_out[4]         = lanes_fifo_response_merge_lane_in_signals_out[4][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[4][0] = lanes_fifo_response_lane_in_signals_in[4];
                      assign lanes_request_lane_out[4]                          = lanes_request_cast_lane_out[4][0];
                      assign lanes_response_merge_engine_in[4][0]               = lanes_response_engine_in[4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[5][0]  = lanes_fifo_request_lane_out_signals_in[5];
                      assign lanes_fifo_request_lane_out_signals_out[5]         = lanes_fifo_request_cast_lane_out_signals_out [5][0];
                      assign lanes_fifo_response_lane_in_signals_out[5]         = lanes_fifo_response_merge_lane_in_signals_out[5][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[5][0] = lanes_fifo_response_lane_in_signals_in[5];
                      assign lanes_request_lane_out[5]                          = lanes_request_cast_lane_out[5][0];
                      assign lanes_response_merge_engine_in[5][0]               = lanes_response_engine_in[5];

                    end
endgenerate

generate
     if(ID_BUNDLE == 1)
                    begin
                      assign lanes_fifo_request_cast_lane_out_signals_in[0][0]  = lanes_fifo_request_lane_out_signals_in[0];
                      assign lanes_fifo_request_lane_out_signals_out[0]         = lanes_fifo_request_cast_lane_out_signals_out [0][0];
                      assign lanes_fifo_response_lane_in_signals_out[0]         = lanes_fifo_response_merge_lane_in_signals_out[0][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][0] = lanes_fifo_response_lane_in_signals_in[0];
                      assign lanes_request_lane_out[0]                          = lanes_request_cast_lane_out[0][0];
                      assign lanes_response_merge_engine_in[0][0]               = lanes_response_engine_in[0];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][2].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][1]                                 = lanes_request_cast_lane_out[1][2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][3].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][2]                                 = lanes_request_cast_lane_out[2][3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][4].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][3].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][3].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][3]                                 = lanes_request_cast_lane_out[3][4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][0]  = lanes_fifo_request_lane_out_signals_in[1];
                      assign lanes_fifo_request_lane_out_signals_out[1]         = lanes_fifo_request_cast_lane_out_signals_out [1][0];
                      assign lanes_fifo_response_lane_in_signals_out[1]         = lanes_fifo_response_merge_lane_in_signals_out[1][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][0] = lanes_fifo_response_lane_in_signals_in[1];
                      assign lanes_request_lane_out[1]                          = lanes_request_cast_lane_out[1][0];
                      assign lanes_response_merge_engine_in[1][0]               = lanes_response_engine_in[1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][4].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][1]                                 = lanes_request_cast_lane_out[2][4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][5].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][2]                                 = lanes_request_cast_lane_out[3][5];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][0]  = lanes_fifo_request_lane_out_signals_in[2];
                      assign lanes_fifo_request_lane_out_signals_out[2]         = lanes_fifo_request_cast_lane_out_signals_out [2][0];
                      assign lanes_fifo_response_lane_in_signals_out[2]         = lanes_fifo_response_merge_lane_in_signals_out[2][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][0] = lanes_fifo_response_lane_in_signals_in[2];
                      assign lanes_request_lane_out[2]                          = lanes_request_cast_lane_out[2][0];
                      assign lanes_response_merge_engine_in[2][0]               = lanes_response_engine_in[2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][6].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[2][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[2][1]                                 = lanes_request_cast_lane_out[3][6];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][0]  = lanes_fifo_request_lane_out_signals_in[3];
                      assign lanes_fifo_request_lane_out_signals_out[3]         = lanes_fifo_request_cast_lane_out_signals_out [3][0];
                      assign lanes_fifo_response_lane_in_signals_out[3]         = lanes_fifo_response_merge_lane_in_signals_out[3][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[3][0] = lanes_fifo_response_lane_in_signals_in[3];
                      assign lanes_request_lane_out[3]                          = lanes_request_cast_lane_out[3][0];
                      assign lanes_response_merge_engine_in[3][0]               = lanes_response_engine_in[3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[4][0]  = lanes_fifo_request_lane_out_signals_in[4];
                      assign lanes_fifo_request_lane_out_signals_out[4]         = lanes_fifo_request_cast_lane_out_signals_out [4][0];
                      assign lanes_fifo_response_lane_in_signals_out[4]         = lanes_fifo_response_merge_lane_in_signals_out[4][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[4][0] = lanes_fifo_response_lane_in_signals_in[4];
                      assign lanes_request_lane_out[4]                          = lanes_request_cast_lane_out[4][0];
                      assign lanes_response_merge_engine_in[4][0]               = lanes_response_engine_in[4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[5][0]  = lanes_fifo_request_lane_out_signals_in[5];
                      assign lanes_fifo_request_lane_out_signals_out[5]         = lanes_fifo_request_cast_lane_out_signals_out [5][0];
                      assign lanes_fifo_response_lane_in_signals_out[5]         = lanes_fifo_response_merge_lane_in_signals_out[5][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[5][0] = lanes_fifo_response_lane_in_signals_in[5];
                      assign lanes_request_lane_out[5]                          = lanes_request_cast_lane_out[5][0];
                      assign lanes_response_merge_engine_in[5][0]               = lanes_response_engine_in[5];

                    end
endgenerate

generate
     if(ID_BUNDLE == 2)
                    begin
                      assign lanes_fifo_request_cast_lane_out_signals_in[0][0]  = lanes_fifo_request_lane_out_signals_in[0];
                      assign lanes_fifo_request_lane_out_signals_out[0]         = lanes_fifo_request_cast_lane_out_signals_out [0][0];
                      assign lanes_fifo_response_lane_in_signals_out[0]         = lanes_fifo_response_merge_lane_in_signals_out[0][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][0] = lanes_fifo_response_lane_in_signals_in[0];
                      assign lanes_request_lane_out[0]                          = lanes_request_cast_lane_out[0][0];
                      assign lanes_response_merge_engine_in[0][0]               = lanes_response_engine_in[0];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][3].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][1]                                 = lanes_request_cast_lane_out[1][3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][5].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][2]                                 = lanes_request_cast_lane_out[2][5];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][7].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][3].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][3].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][3]                                 = lanes_request_cast_lane_out[3][7];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][0]  = lanes_fifo_request_lane_out_signals_in[1];
                      assign lanes_fifo_request_lane_out_signals_out[1]         = lanes_fifo_request_cast_lane_out_signals_out [1][0];
                      assign lanes_fifo_response_lane_in_signals_out[1]         = lanes_fifo_response_merge_lane_in_signals_out[1][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][0] = lanes_fifo_response_lane_in_signals_in[1];
                      assign lanes_request_lane_out[1]                          = lanes_request_cast_lane_out[1][0];
                      assign lanes_response_merge_engine_in[1][0]               = lanes_response_engine_in[1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][6].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][1]                                 = lanes_request_cast_lane_out[2][6];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][8].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][2]                                 = lanes_request_cast_lane_out[3][8];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][0]  = lanes_fifo_request_lane_out_signals_in[2];
                      assign lanes_fifo_request_lane_out_signals_out[2]         = lanes_fifo_request_cast_lane_out_signals_out [2][0];
                      assign lanes_fifo_response_lane_in_signals_out[2]         = lanes_fifo_response_merge_lane_in_signals_out[2][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][0] = lanes_fifo_response_lane_in_signals_in[2];
                      assign lanes_request_lane_out[2]                          = lanes_request_cast_lane_out[2][0];
                      assign lanes_response_merge_engine_in[2][0]               = lanes_response_engine_in[2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][9].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[2][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[2][1]                                 = lanes_request_cast_lane_out[3][9];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][0]  = lanes_fifo_request_lane_out_signals_in[3];
                      assign lanes_fifo_request_lane_out_signals_out[3]         = lanes_fifo_request_cast_lane_out_signals_out [3][0];
                      assign lanes_fifo_response_lane_in_signals_out[3]         = lanes_fifo_response_merge_lane_in_signals_out[3][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[3][0] = lanes_fifo_response_lane_in_signals_in[3];
                      assign lanes_request_lane_out[3]                          = lanes_request_cast_lane_out[3][0];
                      assign lanes_response_merge_engine_in[3][0]               = lanes_response_engine_in[3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[4][0]  = lanes_fifo_request_lane_out_signals_in[4];
                      assign lanes_fifo_request_lane_out_signals_out[4]         = lanes_fifo_request_cast_lane_out_signals_out [4][0];
                      assign lanes_fifo_response_lane_in_signals_out[4]         = lanes_fifo_response_merge_lane_in_signals_out[4][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[4][0] = lanes_fifo_response_lane_in_signals_in[4];
                      assign lanes_request_lane_out[4]                          = lanes_request_cast_lane_out[4][0];
                      assign lanes_response_merge_engine_in[4][0]               = lanes_response_engine_in[4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[5][0]  = lanes_fifo_request_lane_out_signals_in[5];
                      assign lanes_fifo_request_lane_out_signals_out[5]         = lanes_fifo_request_cast_lane_out_signals_out [5][0];
                      assign lanes_fifo_response_lane_in_signals_out[5]         = lanes_fifo_response_merge_lane_in_signals_out[5][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[5][0] = lanes_fifo_response_lane_in_signals_in[5];
                      assign lanes_request_lane_out[5]                          = lanes_request_cast_lane_out[5][0];
                      assign lanes_response_merge_engine_in[5][0]               = lanes_response_engine_in[5];

                    end
endgenerate

generate
     if(ID_BUNDLE == 3)
                    begin
                      assign lanes_fifo_request_cast_lane_out_signals_in[0][0]  = lanes_fifo_request_lane_out_signals_in[0];
                      assign lanes_fifo_request_lane_out_signals_out[0]         = lanes_fifo_request_cast_lane_out_signals_out [0][0];
                      assign lanes_fifo_response_lane_in_signals_out[0]         = lanes_fifo_response_merge_lane_in_signals_out[0][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][0] = lanes_fifo_response_lane_in_signals_in[0];
                      assign lanes_request_lane_out[0]                          = lanes_request_cast_lane_out[0][0];
                      assign lanes_response_merge_engine_in[0][0]               = lanes_response_engine_in[0];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][4].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][1]                                 = lanes_request_cast_lane_out[1][4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][7].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][2]                                 = lanes_request_cast_lane_out[2][7];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][10].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[0][3].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[0][3].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[0][3]                                 = lanes_request_cast_lane_out[3][10];

                      assign lanes_fifo_request_cast_lane_out_signals_in[1][0]  = lanes_fifo_request_lane_out_signals_in[1];
                      assign lanes_fifo_request_lane_out_signals_out[1]         = lanes_fifo_request_cast_lane_out_signals_out [1][0];
                      assign lanes_fifo_response_lane_in_signals_out[1]         = lanes_fifo_response_merge_lane_in_signals_out[1][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][0] = lanes_fifo_response_lane_in_signals_in[1];
                      assign lanes_request_lane_out[1]                          = lanes_request_cast_lane_out[1][0];
                      assign lanes_response_merge_engine_in[1][0]               = lanes_response_engine_in[1];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][8].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][1]                                 = lanes_request_cast_lane_out[2][8];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][11].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[1][2].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[1][2].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[1][2]                                 = lanes_request_cast_lane_out[3][11];

                      assign lanes_fifo_request_cast_lane_out_signals_in[2][0]  = lanes_fifo_request_lane_out_signals_in[2];
                      assign lanes_fifo_request_lane_out_signals_out[2]         = lanes_fifo_request_cast_lane_out_signals_out [2][0];
                      assign lanes_fifo_response_lane_in_signals_out[2]         = lanes_fifo_response_merge_lane_in_signals_out[2][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][0] = lanes_fifo_response_lane_in_signals_in[2];
                      assign lanes_request_lane_out[2]                          = lanes_request_cast_lane_out[2][0];
                      assign lanes_response_merge_engine_in[2][0]               = lanes_response_engine_in[2];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][12].rd_en             = ~lanes_fifo_response_merge_lane_in_signals_out[2][1].prog_full;
                      assign lanes_fifo_response_merge_lane_in_signals_in[2][1].rd_en             = 1'b1;
                      assign lanes_response_merge_engine_in[2][1]                                 = lanes_request_cast_lane_out[3][12];

                      assign lanes_fifo_request_cast_lane_out_signals_in[3][0]  = lanes_fifo_request_lane_out_signals_in[3];
                      assign lanes_fifo_request_lane_out_signals_out[3]         = lanes_fifo_request_cast_lane_out_signals_out [3][0];
                      assign lanes_fifo_response_lane_in_signals_out[3]         = lanes_fifo_response_merge_lane_in_signals_out[3][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[3][0] = lanes_fifo_response_lane_in_signals_in[3];
                      assign lanes_request_lane_out[3]                          = lanes_request_cast_lane_out[3][0];
                      assign lanes_response_merge_engine_in[3][0]               = lanes_response_engine_in[3];

                      assign lanes_fifo_request_cast_lane_out_signals_in[4][0]  = lanes_fifo_request_lane_out_signals_in[4];
                      assign lanes_fifo_request_lane_out_signals_out[4]         = lanes_fifo_request_cast_lane_out_signals_out [4][0];
                      assign lanes_fifo_response_lane_in_signals_out[4]         = lanes_fifo_response_merge_lane_in_signals_out[4][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[4][0] = lanes_fifo_response_lane_in_signals_in[4];
                      assign lanes_request_lane_out[4]                          = lanes_request_cast_lane_out[4][0];
                      assign lanes_response_merge_engine_in[4][0]               = lanes_response_engine_in[4];

                      assign lanes_fifo_request_cast_lane_out_signals_in[5][0]  = lanes_fifo_request_lane_out_signals_in[5];
                      assign lanes_fifo_request_lane_out_signals_out[5]         = lanes_fifo_request_cast_lane_out_signals_out [5][0];
                      assign lanes_fifo_response_lane_in_signals_out[5]         = lanes_fifo_response_merge_lane_in_signals_out[5][0];
                      assign lanes_fifo_response_merge_lane_in_signals_in[5][0] = lanes_fifo_response_lane_in_signals_in[5];
                      assign lanes_request_lane_out[5]                          = lanes_request_cast_lane_out[5][0];
                      assign lanes_response_merge_engine_in[5][0]               = lanes_response_engine_in[5];

                    end
endgenerate
// total_luts=138956

