
        parameter integer C_M00_AXI_ADDR_WIDTH       = 64           ;
        parameter integer C_M00_AXI_DATA_WIDTH       = 512        ;
        parameter integer C_M00_AXI_ID_WIDTH         = M00_AXI4_BE_ID_W          ;
        

        parameter integer C_M01_AXI_ADDR_WIDTH       = 64           ;
        parameter integer C_M01_AXI_DATA_WIDTH       = 512        ;
        parameter integer C_M01_AXI_ID_WIDTH         = M01_AXI4_BE_ID_W          ;
        