
  input  M00_AXI4_MID_MasterReadInterfaceInput   m00_axi_read_in  ,
  output M00_AXI4_MID_MasterReadInterfaceOutput  m00_axi_read_out ,
  input  M00_AXI4_MID_MasterWriteInterfaceInput  m00_axi_write_in ,
  output M00_AXI4_MID_MasterWriteInterfaceOutput m00_axi_write_out,
    

  input  M01_AXI4_MID_MasterReadInterfaceInput   m01_axi_read_in  ,
  output M01_AXI4_MID_MasterReadInterfaceOutput  m01_axi_read_out ,
  input  M01_AXI4_MID_MasterWriteInterfaceInput  m01_axi_write_in ,
  output M01_AXI4_MID_MasterWriteInterfaceOutput m01_axi_write_out,
    