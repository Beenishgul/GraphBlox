// Name ENGINE_FORWARD_DATA ID 14   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 6    mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 15   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 15   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 15   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 1    mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[0][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_READ_WRITE   ID 7    mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[0][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[0][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[0][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[0][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 16   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_READ_WRITE   ID 16   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  1  - Index_Start
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
   // --  2  - Index_End
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  8  - Array_Pointer_RHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_READ_WRITE   ID 16   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_MERGE_DATA   ID 2    mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 8    mapping 4    cycles 2    None-None ( 0 )-( 0 )
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  2  - Index_End
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 3    mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 9    mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 4    mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 10   mapping 2    cycles 10   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[1][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  1  - Index_Start
    graph.overlay_program[1][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[4][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
   // --  2  - Index_End
    graph.overlay_program[1][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[4][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  8  - Array_Pointer_RHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[2][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[4][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[2][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[5][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[5][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
   // --  9  - Array_size
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  2  - Index_End
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
   // --  9  - Array_size
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  9  - Array_size
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 5    mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
   // --  1  - Index_Start
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  2  - Index_End
// Name ENGINE_FILTER_COND  ID 11   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
   // --  9  - Array_size
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 6    mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 12   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 7    mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 13   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[3][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// Name ENGINE_FORWARD_DATA ID 14   mapping 6    cycles 1    None-None ( 0 )-( 0 )
   // --  1  - Index_Start
   // --  1  - Index_Start
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
   // --  2  - Index_End
   // --  2  - Index_End
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
   // --  9  - Array_size
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
   // --  1  - Index_Start
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  2  - Index_End
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_MERGE_DATA   ID 8    mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  7  - Array_Pointer_LHS
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_FILTER_COND  ID 15   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 9    mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 16   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_CSR_INDEX    ID 10   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  1  - Index_Start
   // --  1  - Index_Start
    graph.overlay_program[4][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  2  - Index_End
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[4][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  7  - Array_Pointer_LHS
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[4][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
   // --  8  - Array_Pointer_RHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[5][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
   // --  9  - Array_size
   // --  9  - Array_size
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[5][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 11   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_ALU_OPS      ID 12   mapping 5    cycles 6    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_FILTER_COND  ID 13   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 14   mapping 6    cycles 1    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 15   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
   // --  1  - Index_Start
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  2  - Index_End
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  9  - Array_size
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  9  - Array_size
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  2  - Index_End
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// Name ENGINE_READ_WRITE   ID 16   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  8  - Array_Pointer_RHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  2  - Index_End
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[7][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_MERGE_DATA   ID 17   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 18   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
   // --  2  - Index_End
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
   // --  1  - Index_Start
   // --  9  - Array_size
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  8  - Array_Pointer_RHS
   // --  2  - Index_End
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 19   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[8][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  9  - Array_size
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[9][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
   // --  9  - Array_size
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 20   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 21   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  1  - Index_Start
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
   // --  2  - Index_End
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  8  - Array_Pointer_RHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
   // --  9  - Array_size
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_READ_WRITE   ID 22   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[10][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_MERGE_DATA   ID 23   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
   // --  2  - Index_End
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_FILTER_COND  ID 24   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
   // --  1  - Index_Start
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
   // --  2  - Index_End
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 25   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[11][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[12][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 26   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
   // --  2  - Index_End
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
// Name ENGINE_ALU_OPS      ID 27   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 28   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 29   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 30   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
   // --  2  - Index_End
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
   // --  1  - Index_Start
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
   // --  9  - Array_size
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_READ_WRITE   ID 31   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  2  - Index_End
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  8  - Array_Pointer_RHS
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[14][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  1  - Index_Start
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  2  - Index_End
    graph.overlay_program[15][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 32   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 33   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  2  - Index_End
   // --  8  - Array_Pointer_RHS
   // --  1  - Index_Start
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  9  - Array_size
   // --  2  - Index_End
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
   // --  1  - Index_Start
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  7  - Array_Pointer_LHS
// Name ENGINE_READ_WRITE   ID 34   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  1  - Index_Start
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
   // --  9  - Array_size
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  2  - Index_End
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  9  - Array_size
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[16][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 35   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 36   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
   // --  1  - Index_Start
   // --  2  - Index_End
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
   // --  2  - Index_End
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
   // --  7  - Array_Pointer_LHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
   // --  9  - Array_size
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
   // --  1  - Index_Start
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  2  - Index_End
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
   // --  7  - Array_Pointer_LHS
// Name ENGINE_READ_WRITE   ID 37   mapping 1    cycles 13   None-None ( 0 )-( 0 )
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
   // --  1  - Index_Start
   // --  9  - Array_size
   // --  9  - Array_size
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 );
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*10)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[17][(M_AXI4_FE_DATA_W*15)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*0)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[18][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 38   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// Name ENGINE_FILTER_COND  ID 39   mapping 3    cycles 9    None-None ( 0 )-( 0 )
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
   // --  2  - Index_End
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
   // --  9  - Array_size
   // --  9  - Array_size
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 40   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*1)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*2)+:M_AXI4_FE_DATA_W]  = ( 0 );
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*7)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*8)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[19][(M_AXI4_FE_DATA_W*9)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 41   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// -->  Full  <-- 
   // --  1  - Index_Start
// -->  Full  <-- 
// Number of entries 464
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Number of entries 464
// --------------------------------------------------------------------------------------
   // --  2  - Index_End
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  7  - Array_Pointer_LHS
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  8  - Array_Pointer_RHS
// Name ENGINE_ALU_OPS      ID 42   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
   // --  9  - Array_size
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 43   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 44   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// -->  Full  <-- 
// -->  Full  <-- 
// -->  Full  <-- 
// Number of entries 464
// Number of entries 464
// Number of entries 464
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 45   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 46   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[21][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[22][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 47   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 48   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 49   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[23][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 50   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 51   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_READ_WRITE   ID 52   mapping 1    cycles 13   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[24][(M_AXI4_FE_DATA_W*14)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*3)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*4)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[25][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// -->  Full  <-- 
// Number of entries 464
// --------------------------------------------------------------------------------------
// Name ENGINE_MERGE_DATA   ID 53   mapping 4    cycles 2    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 54   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_CSR_INDEX    ID 55   mapping 2    cycles 10   None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
   // --  1  - Index_Start
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*5)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  2  - Index_End
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*6)+:M_AXI4_FE_DATA_W]  = ( 0 );
   // --  7  - Array_Pointer_LHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*11)+:M_AXI4_FE_DATA_W]  = 0;
   // --  8  - Array_Pointer_RHS
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*12)+:M_AXI4_FE_DATA_W]  = 0;
   // --  9  - Array_size
    graph.overlay_program[26][(M_AXI4_FE_DATA_W*13)+:M_AXI4_FE_DATA_W]  = ( 0 )-( 0 );
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 56   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_ALU_OPS      ID 57   mapping 5    cycles 6    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 58   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FORWARD_DATA ID 59   mapping 6    cycles 1    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// Name ENGINE_FILTER_COND  ID 60   mapping 3    cycles 9    None-None ( 0 )-( 0 )
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
// -->  Full  <-- 
// Number of entries 464
