// -----------------------------------------------------------------------------
//
//      "GLay: A Vertex Centric Re-Configurable Graph Processing Overlay"
//
// -----------------------------------------------------------------------------
// Copyright (c) 2021-2023 All rights reserved
// -----------------------------------------------------------------------------
// Author : Abdullah Mughrabi atmughrabi@gmail.com/atmughra@virginia.edu
// File   : engine_read_write_configure_memory.sv
// Create : 2023-07-17 15:02:02
// Revise : 2023-08-28 15:42:14
// Editor : sublime text4, tab size (4)
// -----------------------------------------------------------------------------

import PKG_AXI4::*;
import PKG_GLOBALS::*;
import PKG_DESCRIPTOR::*;
import PKG_CONTROL::*;
import PKG_MEMORY::*;
import PKG_ENGINE::*;
import PKG_CACHE::*;

module engine_read_write_configure_memory #(parameter
    ID_CU            = 0                                ,
    ID_BUNDLE        = 0                                ,
    ID_LANE          = 0                                ,
    ID_ENGINE        = 0                                ,
    ID_RELATIVE      = 0                                ,
    ID_MODULE        = 0                                ,
    FIFO_WRITE_DEPTH = 16                               ,
    PROG_THRESH      = 8                                ,
    ENGINE_SEQ_WIDTH = 16                               ,
    ENGINE_SEQ_MIN   = ID_RELATIVE * ENGINE_SEQ_WIDTH   ,
    ENGINE_SEQ_MAX   = ENGINE_SEQ_WIDTH + ENGINE_SEQ_MIN
) (
    input  logic                  ap_clk                             ,
    input  logic                  areset                             ,
    input  MemoryPacket           response_memory_in                 ,
    input  FIFOStateSignalsInput  fifo_response_memory_in_signals_in ,
    output FIFOStateSignalsOutput fifo_response_memory_in_signals_out,
    output ReadWriteConfiguration configure_memory_out               ,
    input  FIFOStateSignalsInput  fifo_configure_memory_signals_in   ,
    output FIFOStateSignalsOutput fifo_configure_memory_signals_out  ,
    output logic                  fifo_setup_signal
);

// --------------------------------------------------------------------------------------
// Wires and Variables
// --------------------------------------------------------------------------------------
    logic areset_read_write_generator;
    logic areset_fifo                ;

    MemoryPacket                      response_memory_in_reg                          ;
    MemoryPacketMeta                  configure_memory_meta_int                       ;
    ReadWriteConfiguration            configure_memory_reg                            ;
    ReadWriteConfiguration            configure_memory_int                            ;
    logic [     ENGINE_SEQ_WIDTH-1:0] configure_memory_valid_reg                      ;
    logic [     ENGINE_SEQ_WIDTH-1:0] configure_memory_valid_int                      ;
    logic                             configure_memory_valid_flag                     ;
    logic [CACHE_FRONTEND_ADDR_W-1:0] response_memory_in_reg_offset_sequence          ;
    logic [CACHE_FRONTEND_ADDR_W-1:0] fifo_response_memory_in_dout_int_offset_sequence;

// --------------------------------------------------------------------------------------
// Response FIFO
// --------------------------------------------------------------------------------------
    MemoryPacketPayload    fifo_response_memory_in_din             ;
    MemoryPacket           fifo_response_memory_in_dout_int        ;
    MemoryPacketPayload    fifo_response_memory_in_dout            ;
    FIFOStateSignalsInput  fifo_response_memory_in_signals_in_reg  ;
    FIFOStateSignalsInput  fifo_response_memory_in_signals_in_int  ;
    FIFOStateSignalsOutput fifo_response_memory_in_signals_out_int ;
    logic                  fifo_response_memory_in_setup_signal_int;
    logic                  fifo_response_memory_in_push_filter     ;

// --------------------------------------------------------------------------------------
// Configure FIFO
// --------------------------------------------------------------------------------------
    ReadWriteConfigurationPayload fifo_configure_memory_din             ;
    ReadWriteConfiguration        fifo_configure_memory_dout_int        ;
    ReadWriteConfigurationPayload fifo_configure_memory_dout            ;
    FIFOStateSignalsInput         fifo_configure_memory_signals_in_reg  ;
    FIFOStateSignalsInput         fifo_configure_memory_signals_in_int  ;
    FIFOStateSignalsOutput        fifo_configure_memory_signals_out_int ;
    logic                         fifo_configure_memory_setup_signal_int;

// --------------------------------------------------------------------------------------
// Register reset signal
// --------------------------------------------------------------------------------------
    always_ff @(posedge ap_clk) begin
        areset_read_write_generator <= areset;
        areset_fifo                 <= areset;
    end

// --------------------------------------------------------------------------------------
// Drive input
// --------------------------------------------------------------------------------------
    always_ff @(posedge ap_clk) begin
        if(areset_read_write_generator) begin
            response_memory_in_reg.valid           <= 1'b0;
            fifo_response_memory_in_signals_in_reg <= 0;
            fifo_configure_memory_signals_in_reg   <= 0;
        end else begin
            response_memory_in_reg.valid                 <= response_memory_in.valid ;
            fifo_response_memory_in_signals_in_reg.rd_en <= fifo_response_memory_in_signals_in.rd_en;
            fifo_configure_memory_signals_in_reg.rd_en   <= fifo_configure_memory_signals_in.rd_en;
        end
    end

    always_ff @(posedge ap_clk) begin
        response_memory_in_reg.payload <= response_memory_in.payload;
    end

// --------------------------------------------------------------------------------------
// Drive output
// --------------------------------------------------------------------------------------
    always_ff @(posedge ap_clk) begin
        if(areset_read_write_generator) begin
            fifo_setup_signal          <= 1'b1;
            configure_memory_out.valid <= 0;
        end else begin
            fifo_setup_signal          <= fifo_response_memory_in_setup_signal_int | fifo_configure_memory_setup_signal_int;
            configure_memory_out.valid <= fifo_configure_memory_dout_int.valid;
        end
    end

    always_ff @(posedge ap_clk) begin
        fifo_response_memory_in_signals_out <= fifo_response_memory_in_signals_out_int;
        fifo_configure_memory_signals_out   <= fifo_configure_memory_signals_out_int;
        configure_memory_out.payload        <= fifo_configure_memory_dout_int.payload;
    end


// --------------------------------------------------------------------------------------
// Create Configuration Packet
// --------------------------------------------------------------------------------------
    assign configure_memory_valid_flag                      = &configure_memory_valid_reg;
    assign response_memory_in_reg_offset_sequence           = (response_memory_in_reg.payload.meta.address.offset >> response_memory_in_reg.payload.meta.address.shift.amount);
    assign fifo_response_memory_in_dout_int_offset_sequence = (fifo_response_memory_in_dout_int.payload.meta.address.offset >> fifo_response_memory_in_dout_int.payload.meta.address.shift.amount);

    always_comb begin
        configure_memory_meta_int.route.from.id_cu        = 1'b1 << ID_CU;
        configure_memory_meta_int.route.from.id_bundle    = 1'b1 << ID_BUNDLE;
        configure_memory_meta_int.route.from.id_lane      = 1'b1 << ID_LANE;
        configure_memory_meta_int.route.from.id_engine    = 1'b1 << ID_ENGINE;
        configure_memory_meta_int.route.from.id_module    = 1'b1 << ID_MODULE;
        configure_memory_meta_int.route.from.id_buffer    = 0;
        configure_memory_meta_int.route.to.id_cu          = 0;
        configure_memory_meta_int.route.to.id_bundle      = 0;
        configure_memory_meta_int.route.to.id_lane        = 0;
        configure_memory_meta_int.route.to.id_engine      = 0;
        configure_memory_meta_int.route.to.id_module      = 1;
        configure_memory_meta_int.route.to.id_buffer      = 0;
        configure_memory_meta_int.route.seq_src.id_cu     = 1'b1 << ID_CU;
        configure_memory_meta_int.route.seq_src.id_bundle = 1'b1 << ID_BUNDLE;
        configure_memory_meta_int.route.seq_src.id_lane   = 1'b1 << ID_LANE;
        configure_memory_meta_int.route.seq_src.id_engine = 1'b1 << ID_ENGINE;
        configure_memory_meta_int.route.seq_src.id_module = 1'b1 << ID_MODULE;
        configure_memory_meta_int.route.seq_src.id_buffer = 0;
        configure_memory_meta_int.route.seq_state         = SEQUENCE_INVALID;
        configure_memory_meta_int.route.hops              = CU_BUNDLE_COUNT_WIDTH_BITS;
        configure_memory_meta_int.address.base            = 0;
        configure_memory_meta_int.address.offset          = $clog2(CACHE_FRONTEND_DATA_W/8);
        configure_memory_meta_int.address.shift.amount    = 0;
        configure_memory_meta_int.address.shift.direction = 1'b1;
        configure_memory_meta_int.subclass.cmd            = CMD_INVALID;
        configure_memory_meta_int.subclass.buffer         = STRUCT_INVALID;
    end

    always_comb begin
        configure_memory_int.valid                        = configure_memory_valid_int;
        configure_memory_int.payload.meta.route.from      = configure_memory_meta_int.route.from;
        configure_memory_int.payload.meta.route.seq_src   = configure_memory_meta_int.route.seq_src;
        configure_memory_int.payload.meta.route.seq_state = configure_memory_meta_int.route.seq_state;
        configure_memory_int.payload.meta.route.hops      = configure_memory_meta_int.route.hops;
        configure_memory_int.payload.meta.address.base    = configure_memory_meta_int.address.base;
        configure_memory_int.payload.meta.address.offset  = configure_memory_meta_int.address.offset;

        if(fifo_response_memory_in_dout_int.valid) begin
            case (fifo_response_memory_in_dout_int_offset_sequence)
                (ENGINE_SEQ_MIN+0) : begin
                    configure_memory_int.payload.param.increment     = fifo_response_memory_in_dout_int.payload.data.field[0][0];
                    configure_memory_int.payload.param.decrement     = fifo_response_memory_in_dout_int.payload.data.field[0][1];
                    configure_memory_int.payload.param.mode_sequence = fifo_response_memory_in_dout_int.payload.data.field[0][2];
                    configure_memory_int.payload.param.mode_buffer   = fifo_response_memory_in_dout_int.payload.data.field[0][3];
                    configure_memory_valid_int[0]                    = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+1) : begin
                    configure_memory_int.payload.param.index_start = fifo_response_memory_in_dout_int.payload.data.field[0];
                    configure_memory_valid_int[1]                  = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+2) : begin
                    configure_memory_int.payload.param.index_end = fifo_response_memory_in_dout_int.payload.data.field[0];
                    configure_memory_valid_int[2]                = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+3) : begin
                    configure_memory_int.payload.param.stride = fifo_response_memory_in_dout_int.payload.data.field[0];
                    configure_memory_valid_int[3]             = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+4) : begin
                    configure_memory_int.payload.param.granularity            = fifo_response_memory_in_dout_int.payload.data.field[0][CACHE_FRONTEND_DATA_W-2:0];
                    configure_memory_int.payload.meta.address.shift.amount    = fifo_response_memory_in_dout_int.payload.data.field[0][CACHE_FRONTEND_DATA_W-2:0];
                    configure_memory_int.payload.meta.address.shift.direction = fifo_response_memory_in_dout_int.payload.data.field[0][CACHE_FRONTEND_DATA_W-1];
                    configure_memory_valid_int[4]                             = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+5) : begin
                    configure_memory_int.payload.meta.subclass.cmd    = type_memory_cmd'(fifo_response_memory_in_dout_int.payload.data.field[0][TYPE_MEMORY_CMD_BITS-1:0]);
                    configure_memory_int.payload.meta.subclass.buffer = type_data_buffer'(fifo_response_memory_in_dout_int.payload.data.field[0][(TYPE_DATA_STRUCTURE_BITS+TYPE_MEMORY_CMD_BITS)-1:TYPE_MEMORY_CMD_BITS]);
                    configure_memory_valid_int[5]                     = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+6) : begin
                    configure_memory_valid_int[6] = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+7) : begin
                    configure_memory_int.payload.meta.route.to.id_cu     = fifo_response_memory_in_dout_int.payload.data.field[0][(CU_KERNEL_COUNT_WIDTH_BITS)-1:0];
                    configure_memory_int.payload.meta.route.to.id_bundle = fifo_response_memory_in_dout_int.payload.data.field[0][(CU_BUNDLE_COUNT_WIDTH_BITS+CU_KERNEL_COUNT_WIDTH_BITS)-1:CU_KERNEL_COUNT_WIDTH_BITS];
                    configure_memory_int.payload.meta.route.to.id_lane   = fifo_response_memory_in_dout_int.payload.data.field[0][(CU_LANE_COUNT_WIDTH_BITS+CU_BUNDLE_COUNT_WIDTH_BITS+CU_KERNEL_COUNT_WIDTH_BITS)-1:(CU_BUNDLE_COUNT_WIDTH_BITS+CU_KERNEL_COUNT_WIDTH_BITS)];
                    configure_memory_int.payload.meta.route.to.id_buffer = fifo_response_memory_in_dout_int.payload.data.field[0][(CU_BUFFER_COUNT_WIDTH_BITS+CU_LANE_COUNT_WIDTH_BITS+CU_BUNDLE_COUNT_WIDTH_BITS+CU_KERNEL_COUNT_WIDTH_BITS)-1:(CU_LANE_COUNT_WIDTH_BITS+CU_BUNDLE_COUNT_WIDTH_BITS+CU_KERNEL_COUNT_WIDTH_BITS)];
                    configure_memory_valid_int[7]                        = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+8) : begin
                    configure_memory_int.payload.param.array_pointer[(CACHE_FRONTEND_DATA_W)-1:0] = fifo_response_memory_in_dout_int.payload.data.field[0];
                    configure_memory_valid_int[8]                                                 = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+9) : begin
                    configure_memory_int.payload.param.array_pointer[(M_AXI_MEMORY_ADDR_WIDTH)-1:CACHE_FRONTEND_DATA_W] = fifo_response_memory_in_dout_int.payload.data.field[0];
                    configure_memory_valid_int[9]                                                                       = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+10) : begin
                    configure_memory_int.payload.param.array_size = fifo_response_memory_in_dout_int.payload.data.field[0];
                    configure_memory_valid_int[10]                = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+11) : begin
                    configure_memory_valid_int[11] = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+12) : begin
                    configure_memory_valid_int[12] = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+13) : begin
                    configure_memory_valid_int[13] = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+14) : begin
                    configure_memory_valid_int[14] = 1'b1  ;
                end
                (ENGINE_SEQ_MIN+15) : begin
                    configure_memory_valid_int[15] = 1'b1  ;
                end
                default : begin
                    configure_memory_int.payload.param = configure_memory_int.payload.param;
                    if(configure_memory_valid_int)
                        configure_memory_valid_int = 0;
                    else
                        configure_memory_valid_int = configure_memory_valid_int;
                end
            endcase
        end else begin
            configure_memory_int.payload.param = configure_memory_int.payload.param;
            if(configure_memory_valid_int)
                configure_memory_valid_int = 0;
            else
                configure_memory_valid_int = configure_memory_valid_int;
        end
    end

    always_ff @(posedge ap_clk) begin
        if(areset_read_write_generator) begin
            configure_memory_valid_reg <= 0;
            configure_memory_reg.valid <= 1'b0;
        end else begin
            configure_memory_valid_reg <= configure_memory_valid_int;
            configure_memory_reg.valid <= configure_memory_int.valid;
        end
    end

    always_ff @(posedge ap_clk) begin
        configure_memory_reg.payload <= configure_memory_int.payload;
    end

// --------------------------------------------------------------------------------------
// FIFO memory response out fifo MemoryPacket
// --------------------------------------------------------------------------------------
    // FIFO is resetting
    assign fifo_response_memory_in_setup_signal_int = fifo_response_memory_in_signals_out_int.wr_rst_busy  | fifo_response_memory_in_signals_out_int.rd_rst_busy;

    // Push
    assign fifo_response_memory_in_push_filter          = ((response_memory_in_reg.payload.meta.subclass.buffer == STRUCT_CU_SETUP)|(response_memory_in_reg.payload.meta.subclass.buffer == STRUCT_ENGINE_SETUP)) & (response_memory_in_reg_offset_sequence < (ENGINE_SEQ_MAX)) & (response_memory_in_reg_offset_sequence >= ENGINE_SEQ_MIN);
    assign fifo_response_memory_in_signals_in_int.wr_en = response_memory_in_reg.valid & fifo_response_memory_in_push_filter;
    assign fifo_response_memory_in_din                  = response_memory_in_reg.payload;

    // Pop
    assign fifo_response_memory_in_signals_in_int.rd_en = ~fifo_response_memory_in_signals_out_int.empty & fifo_response_memory_in_signals_in_reg.rd_en & ~(configure_memory_valid_flag) & ~fifo_configure_memory_signals_out_int.prog_full ;
    assign fifo_response_memory_in_dout_int.valid       = fifo_response_memory_in_signals_out_int.valid;
    assign fifo_response_memory_in_dout_int.payload     = fifo_response_memory_in_dout;

    xpm_fifo_sync_wrapper #(
        .FIFO_WRITE_DEPTH(FIFO_WRITE_DEPTH          ),
        .WRITE_DATA_WIDTH($bits(MemoryPacketPayload)),
        .READ_DATA_WIDTH ($bits(MemoryPacketPayload)),
        .PROG_THRESH     (PROG_THRESH               )
    ) inst_fifo_MemoryPacketResponseMemoryInput (
        .clk        (ap_clk                                             ),
        .srst       (areset_fifo                                        ),
        .din        (fifo_response_memory_in_din                        ),
        .wr_en      (fifo_response_memory_in_signals_in_int.wr_en       ),
        .rd_en      (fifo_response_memory_in_signals_in_int.rd_en       ),
        .dout       (fifo_response_memory_in_dout                       ),
        .full       (fifo_response_memory_in_signals_out_int.full       ),
        .empty      (fifo_response_memory_in_signals_out_int.empty      ),
        .valid      (fifo_response_memory_in_signals_out_int.valid      ),
        .prog_full  (fifo_response_memory_in_signals_out_int.prog_full  ),
        .wr_rst_busy(fifo_response_memory_in_signals_out_int.wr_rst_busy),
        .rd_rst_busy(fifo_response_memory_in_signals_out_int.rd_rst_busy)
    );

// --------------------------------------------------------------------------------------
// FIFO memory configure_memory out fifo MemoryPacket
// --------------------------------------------------------------------------------------
    // FIFO is resetting
    assign fifo_configure_memory_setup_signal_int = fifo_configure_memory_signals_out_int.wr_rst_busy  | fifo_configure_memory_signals_out_int.rd_rst_busy;

    // Push
    assign fifo_configure_memory_signals_in_int.wr_en = configure_memory_reg.valid;
    assign fifo_configure_memory_din                  = configure_memory_reg.payload;

    // Pop
    assign fifo_configure_memory_signals_in_int.rd_en = ~fifo_configure_memory_signals_out_int.empty & fifo_configure_memory_signals_in_reg.rd_en;
    assign fifo_configure_memory_dout_int.valid       = fifo_configure_memory_signals_out_int.valid;
    assign fifo_configure_memory_dout_int.payload     = fifo_configure_memory_dout;

    xpm_fifo_sync_wrapper #(
        .FIFO_WRITE_DEPTH(FIFO_WRITE_DEPTH                    ),
        .WRITE_DATA_WIDTH($bits(ReadWriteConfigurationPayload)),
        .READ_DATA_WIDTH ($bits(ReadWriteConfigurationPayload)),
        .PROG_THRESH     (PROG_THRESH                         )
    ) inst_fifo_MemoryPacketResponseConigurationInput (
        .clk        (ap_clk                                           ),
        .srst       (areset_fifo                                      ),
        .din        (fifo_configure_memory_din                        ),
        .wr_en      (fifo_configure_memory_signals_in_int.wr_en       ),
        .rd_en      (fifo_configure_memory_signals_in_int.rd_en       ),
        .dout       (fifo_configure_memory_dout                       ),
        .full       (fifo_configure_memory_signals_out_int.full       ),
        .empty      (fifo_configure_memory_signals_out_int.empty      ),
        .valid      (fifo_configure_memory_signals_out_int.valid      ),
        .prog_full  (fifo_configure_memory_signals_out_int.prog_full  ),
        .wr_rst_busy(fifo_configure_memory_signals_out_int.wr_rst_busy),
        .rd_rst_busy(fifo_configure_memory_signals_out_int.rd_rst_busy)
    );

endmodule : engine_read_write_configure_memory