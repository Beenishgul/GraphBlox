// -----------------------------------------------------------------------------
//
//      "GLay: A Vertex Centric Re-Configurable Graph Processing Overlay"
//
// -----------------------------------------------------------------------------
// Copyright (c) 2021-2023 All rights reserved
// -----------------------------------------------------------------------------
// Author : Abdullah Mughrabi atmughrabi@gmail.com/atmughra@virginia.edu
// File   : 01_pkg_globals.sv
// Create : 2022-11-16 19:43:34
// Revise : 2023-08-28 14:41:10
// Editor : sublime text4, tab size (4)
// -----------------------------------------------------------------------------
package PKG_GLOBALS;

// ********************************************************************************************
// ***************                  GLOBAL MEMORY(DDR4/HBM)                      **************
// ***************                  ALVEO 250 -> 4  banks (300MHz)               **************
// ***************                  ALVEO 280 -> 32 banks (300/500MHz)           **************
// ********************************************************************************************

// --------------------------------------------------------------------------------------
//  COMPUTE UNITS GLOBALS
// --------------------------------------------------------------------------------------
// Kernel current settings engines/lanes/bundles/buffers
// --------------------------------------------------------------------------------------
	parameter KERNEL_CU_COUNT = 1 ;
	parameter CU_BUNDLE_COUNT = 4 ;
	parameter CU_ENGINE_COUNT = 8 ;
	parameter CU_BUFFER_COUNT = 10;

// --------------------------------------------------------------------------------------
// Maximum supported engines/lanes/bundles/buffers
// --------------------------------------------------------------------------------------
	parameter CU_KERNEL_COUNT_TOTAL       = 8 ;
	parameter CU_BUNDLE_COUNT_TOTAL       = 8 ;
	parameter CU_LANE_COUNT_TOTAL         = 8 ;
	parameter CU_ENGINE_COUNT_TOTAL       = 8 ;
	parameter CU_MODULE_COUNT_TOTAL       = 8 ;
	parameter CU_BUFFER_COUNT_TOTAL       = 8 ;
	parameter CU_PACKET_SEQ_ID_WIDTH_BITS = 16;

// --------------------------------------------------------------------------------------
	parameter CU_KERNEL_COUNT_WIDTH_BITS = CU_KERNEL_COUNT_TOTAL;
	parameter CU_BUNDLE_COUNT_WIDTH_BITS = CU_BUNDLE_COUNT_TOTAL;
	parameter CU_LANE_COUNT_WIDTH_BITS   = CU_LANE_COUNT_TOTAL  ;
	parameter CU_ENGINE_COUNT_WIDTH_BITS = CU_ENGINE_COUNT_TOTAL;
	parameter CU_MODULE_COUNT_WIDTH_BITS = CU_MODULE_COUNT_TOTAL;
	parameter CU_BUFFER_COUNT_WIDTH_BITS = CU_BUFFER_COUNT_TOTAL;

// --------------------------------------------------------------------------------------
//  KERNEL COMMON GLOBALS
// --------------------------------------------------------------------------------------
//  CU -> Cache Changing these values would change the cache front end
// --------------------------------------------------------------------------------------
	parameter GLOBAL_SYSTEM_CACHE_IP = 1 ;
	parameter GLOBAL_CU_CACHE_IP     = 1 ;
// --------------------------------------------------------------------------------------

endpackage