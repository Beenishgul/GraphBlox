.ID_CU                               (ID_CU                               ),
.ID_BUNDLE                           (ID_BUNDLE                           ),
.ID_LANE                             (i                                   ),
.NUM_BUNDLES                         (NUM_BUNDLES                         ),
.NUM_LANES                           (NUM_LANES                           ),
.NUM_ENGINES                         (ENGINES_COUNT_ARRAY[i]              ),
.LANES_COUNT_ARRAY                   (LANES_COUNT_ARRAY                   ),
.ENGINES_COUNT_ARRAY                 (ENGINES_COUNT_ARRAY                 ),
.LANES_ENGINES_COUNT_ARRAY           (LANES_ENGINES_COUNT_ARRAY           ),
.ENGINES_CONFIG_ARRAY                (LANES_CONFIG_ARRAY[i]               ),
.ENGINES_ENGINE_ID_ARRAY             (LANES_ENGINE_ID_ARRAY[i]            ),
.LANES_CONFIG_ARRAY                  (LANES_CONFIG_ARRAY                  ),
.LANES_ENGINE_ID_ARRAY               (LANES_ENGINE_ID_ARRAY               ),
.BUNDLES_CONFIG_ARRAY                (BUNDLES_CONFIG_ARRAY                ),
.BUNDLES_ENGINE_ID_ARRAY             (BUNDLES_ENGINE_ID_ARRAY             ),
.CU_BUNDLES_COUNT_ARRAY              (CU_BUNDLES_COUNT_ARRAY              ),
.CU_BUNDLES_LANES_COUNT_ARRAY        (CU_BUNDLES_LANES_COUNT_ARRAY        ),
.CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY(CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY),
.CU_BUNDLES_CONFIG_ARRAY             (CU_BUNDLES_CONFIG_ARRAY             ),
.CU_BUNDLES_ENGINE_ID_ARRAY          (CU_BUNDLES_ENGINE_ID_ARRAY          )