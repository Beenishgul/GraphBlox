    parameter ID_CU     = 0,
    parameter ID_BUNDLE = 0,
// --------------------------------------------------------------------------------------
// CU SETTINGS
// --------------------------------------------------------------------------------------
`include "topology_parameters.vh"

