.CU_BUNDLES_CONFIG_ARRAY                 (CU_BUNDLES_CONFIG_ARRAY                          ),
.CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN  (CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN           ),       
.CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH(CU_BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH         ),  
.CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST (CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST ),
.CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE(CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE),
.CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE (CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE  ),
.CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY (CU_BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY  ),
.CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE (CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE  ),
.CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY (CU_BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY  ),
.CU_BUNDLES_CONFIG_CAST_WIDTH_ARRAY      (CU_BUNDLES_CONFIG_CAST_WIDTH_ARRAY               ),
.CU_BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST  (CU_BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST ),
.CU_BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE (CU_BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE),
.CU_BUNDLES_CONFIG_CU_ARBITER_NUM_ENGINE     (CU_BUNDLES_CONFIG_CU_ARBITER_NUM_ENGINE      ),
.CU_BUNDLES_CONFIG_CU_ARBITER_NUM_MEMORY     (CU_BUNDLES_CONFIG_CU_ARBITER_NUM_MEMORY      ),
.CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST  (CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE (CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE     (CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE      ),
.CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY     (CU_BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY      ),
.CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST (CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST ),
.CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE(CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE),
.CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_ENGINE (CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_ENGINE  ),
.CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_MEMORY (CU_BUNDLES_CONFIG_ENGINE_ARBITER_NUM_MEMORY  ),
.CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE (CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE  ),
.CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY (CU_BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY  ),
.CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST  (CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST   ),
.CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE  (CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE   ),
.CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_ENGINE   (CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_ENGINE    ),
.CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_MEMORY   (CU_BUNDLES_CONFIG_LANE_ARBITER_NUM_MEMORY    ),
.CU_BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY (CU_BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY          ),
.CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST  (CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST   ),
.CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE  (CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE   ),
.CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE   (CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE    ),
.CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY   (CU_BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY    ),
.CU_BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY  (CU_BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY ),
.CU_BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY (CU_BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY),
.CU_BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY(CU_BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY         ),
.CU_BUNDLES_CONFIG_MAX_CAST_WIDTH_ARRAY  (CU_BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY          ),
.CU_BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY (CU_BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY          ),
.CU_BUNDLES_CONFIG_MERGE_CONNECT_ARRAY   (CU_BUNDLES_CONFIG_MERGE_CONNECT_ARRAY            ),
.CU_BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY (CU_BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY),
.CU_BUNDLES_CONFIG_MERGE_WIDTH_ARRAY     (CU_BUNDLES_CONFIG_MERGE_WIDTH_ARRAY              ),
.CU_BUNDLES_COUNT_ARRAY                  (CU_BUNDLES_COUNT_ARRAY                           ),
.CU_BUNDLES_ENGINE_ID_ARRAY              (CU_BUNDLES_ENGINE_ID_ARRAY                       ),
.CU_BUNDLES_LANES_COUNT_ARRAY            (CU_BUNDLES_LANES_COUNT_ARRAY                     ),
.CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY    (CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY             ),
.BUNDLES_CONFIG_ARRAY                    (BUNDLES_CONFIG_ARRAY                             ),
.BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN     (BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_MIN              ),        
.BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH   (BUNDLES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH            ), 
.BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST (BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST ),
.BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE(BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE ),
.BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE (BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE  ),
.BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY (BUNDLES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY  ),
.BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE ),
.BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE (BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE  ),
.BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY (BUNDLES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY  ),
.BUNDLES_CONFIG_CAST_WIDTH_ARRAY         (BUNDLES_CONFIG_CAST_WIDTH_ARRAY                  ),
.BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST    (BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST  ),
.BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE   (BUNDLES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE ),
.BUNDLES_CONFIG_CU_ARBITER_NUM_ENGINE     (BUNDLES_CONFIG_CU_ARBITER_NUM_ENGINE      ),
.BUNDLES_CONFIG_CU_ARBITER_NUM_MEMORY     (BUNDLES_CONFIG_CU_ARBITER_NUM_MEMORY      ),
.BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST    (BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST  ),
.BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE   (BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE ),
.BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE     (BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE      ),
.BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY     (BUNDLES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY      ),
.BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST (BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST ),
.BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE(BUNDLES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE),
.BUNDLES_CONFIG_ENGINE_ARBITER_NUM_ENGINE (BUNDLES_CONFIG_ENGINE_ARBITER_NUM_ENGINE  ),
.BUNDLES_CONFIG_ENGINE_ARBITER_NUM_MEMORY (BUNDLES_CONFIG_ENGINE_ARBITER_NUM_MEMORY  ),
.BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE (BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE  ),
.BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY (BUNDLES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY  ),
.BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST  (BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST   ),
.BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE  (BUNDLES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE   ),
.BUNDLES_CONFIG_LANE_ARBITER_NUM_ENGINE   (BUNDLES_CONFIG_LANE_ARBITER_NUM_ENGINE    ),
.BUNDLES_CONFIG_LANE_ARBITER_NUM_MEMORY   (BUNDLES_CONFIG_LANE_ARBITER_NUM_MEMORY    ),
.BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY    (BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY             ),
.BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST  (BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST   ),
.BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE  (BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE   ),
.BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE   (BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE    ),
.BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY   (BUNDLES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY    ),
.BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY  (BUNDLES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY       ),
.BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY (BUNDLES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY      ),
.BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY   (BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY            ),
.BUNDLES_CONFIG_MAX_CAST_WIDTH_ARRAY     (BUNDLES_CONFIG_MAX_CAST_WIDTH_ARRAY              ),
.BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY    (BUNDLES_CONFIG_MAX_MERGE_WIDTH_ARRAY             ),
.BUNDLES_CONFIG_MERGE_CONNECT_ARRAY      (BUNDLES_CONFIG_MERGE_CONNECT_ARRAY               ),
.BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY (BUNDLES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY      ),
.BUNDLES_CONFIG_MERGE_WIDTH_ARRAY        (BUNDLES_CONFIG_MERGE_WIDTH_ARRAY                 ),
.BUNDLES_ENGINE_ID_ARRAY                 (BUNDLES_ENGINE_ID_ARRAY                          ),
.LANES_CONFIG_ARRAY                      (LANES_CONFIG_ARRAY                               ),
.LANES_CONFIG_ARRAY_ENGINE_SEQ_MIN       (LANES_CONFIG_ARRAY_ENGINE_SEQ_MIN                ),             
.LANES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH     (LANES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH              ),  
.LANES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST (LANES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST ),
.LANES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE(LANES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE),
.LANES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE (LANES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE  ),
.LANES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY (LANES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY  ),
.LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE (LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE  ),
.LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY (LANES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY  ),
.LANES_CONFIG_CAST_WIDTH_ARRAY           (LANES_CONFIG_CAST_WIDTH_ARRAY                    ),
.LANES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST    (LANES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST  ),
.LANES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE    (LANES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE),
.LANES_CONFIG_CU_ARBITER_NUM_ENGINE     (LANES_CONFIG_CU_ARBITER_NUM_ENGINE      ),
.LANES_CONFIG_CU_ARBITER_NUM_MEMORY     (LANES_CONFIG_CU_ARBITER_NUM_MEMORY      ),
.LANES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST    (LANES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST  ),
.LANES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE    (LANES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.LANES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE     (LANES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE      ),
.LANES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY     (LANES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY      ),
.LANES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST (LANES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST ),
.LANES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE(LANES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE),
.LANES_CONFIG_ENGINE_ARBITER_NUM_ENGINE (LANES_CONFIG_ENGINE_ARBITER_NUM_ENGINE  ),
.LANES_CONFIG_ENGINE_ARBITER_NUM_MEMORY (LANES_CONFIG_ENGINE_ARBITER_NUM_MEMORY  ),
.LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE (LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE  ),
.LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY (LANES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY  ),
.LANES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST  (LANES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST   ),
.LANES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE  (LANES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE   ),
.LANES_CONFIG_LANE_ARBITER_NUM_ENGINE   (LANES_CONFIG_LANE_ARBITER_NUM_ENGINE    ),
.LANES_CONFIG_LANE_ARBITER_NUM_MEMORY   (LANES_CONFIG_LANE_ARBITER_NUM_MEMORY    ),
.LANES_CONFIG_LANE_CAST_WIDTH_ARRAY      (LANES_CONFIG_LANE_CAST_WIDTH_ARRAY               ),
.LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST  (LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST   ),
.LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE  (LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE   ),
.LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE   (LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE    ),
.LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY   (LANES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY    ),
.LANES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY  (LANES_CONFIG_LANE_MAX_CAST_WIDTH_ARRAY           ),
.LANES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY (LANES_CONFIG_LANE_MAX_MERGE_WIDTH_ARRAY          ),
.LANES_CONFIG_LANE_MERGE_WIDTH_ARRAY     (LANES_CONFIG_LANE_MERGE_WIDTH_ARRAY              ),
.LANES_CONFIG_MAX_CAST_WIDTH_ARRAY       (LANES_CONFIG_MAX_CAST_WIDTH_ARRAY                ),
.LANES_CONFIG_MAX_MERGE_WIDTH_ARRAY      (LANES_CONFIG_MAX_MERGE_WIDTH_ARRAY               ),
.LANES_CONFIG_MERGE_CONNECT_ARRAY        (LANES_CONFIG_MERGE_CONNECT_ARRAY                 ),
.LANES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY (LANES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY          ),
.LANES_CONFIG_MERGE_WIDTH_ARRAY          (LANES_CONFIG_MERGE_WIDTH_ARRAY                   ),
.LANES_COUNT_ARRAY                       (LANES_COUNT_ARRAY                                ),
.LANES_ENGINE_ID_ARRAY                   (LANES_ENGINE_ID_ARRAY                            ),
.LANES_ENGINES_COUNT_ARRAY               (LANES_ENGINES_COUNT_ARRAY                        ),
.ENGINES_CONFIG_ARRAY                    (ENGINES_CONFIG_ARRAY                             ),
.ENGINES_CONFIG_ARRAY_ENGINE_SEQ_MIN     (ENGINES_CONFIG_ARRAY_ENGINE_SEQ_MIN              ),                      
.ENGINES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH   (ENGINES_CONFIG_ARRAY_ENGINE_SEQ_WIDTH            ),   
.ENGINES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST (ENGINES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_REQUEST ),
.ENGINES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE(ENGINES_CONFIG_BUNDLE_ARBITER_NUM_CONTROL_RESPONSE),
.ENGINES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE (ENGINES_CONFIG_BUNDLE_ARBITER_NUM_ENGINE  ),
.ENGINES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY (ENGINES_CONFIG_BUNDLE_ARBITER_NUM_MEMORY  ),
.ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE (ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_ENGINE  ),
.ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY (ENGINES_CONFIG_BUNDLE_FIFO_ARBITER_SIZE_MEMORY  ),
.ENGINES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST    (ENGINES_CONFIG_CU_ARBITER_NUM_CONTROL_REQUEST  ),
.ENGINES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE    (ENGINES_CONFIG_CU_ARBITER_NUM_CONTROL_RESPONSE),
.ENGINES_CONFIG_CU_ARBITER_NUM_ENGINE     (ENGINES_CONFIG_CU_ARBITER_NUM_ENGINE      ),
.ENGINES_CONFIG_CU_ARBITER_NUM_MEMORY     (ENGINES_CONFIG_CU_ARBITER_NUM_MEMORY      ),
.ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST    (ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_REQUEST  ),
.ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE    (ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE     (ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_ENGINE      ),
.ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY     (ENGINES_CONFIG_CU_FIFO_ARBITER_SIZE_MEMORY      ),
.ENGINES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST (ENGINES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_REQUEST ),
.ENGINES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE(ENGINES_CONFIG_ENGINE_ARBITER_NUM_CONTROL_RESPONSE),
.ENGINES_CONFIG_ENGINE_ARBITER_NUM_ENGINE (ENGINES_CONFIG_ENGINE_ARBITER_NUM_ENGINE  ),
.ENGINES_CONFIG_ENGINE_ARBITER_NUM_MEMORY (ENGINES_CONFIG_ENGINE_ARBITER_NUM_MEMORY  ),
.ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST (ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_REQUEST ),
.ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE(ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE),
.ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE (ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_ENGINE  ),
.ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY (ENGINES_CONFIG_ENGINE_FIFO_ARBITER_SIZE_MEMORY  ),
.ENGINES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST  (ENGINES_CONFIG_LANE_ARBITER_NUM_CONTROL_REQUEST   ),
.ENGINES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE  (ENGINES_CONFIG_LANE_ARBITER_NUM_CONTROL_RESPONSE ),
.ENGINES_CONFIG_LANE_ARBITER_NUM_ENGINE   (ENGINES_CONFIG_LANE_ARBITER_NUM_ENGINE    ),
.ENGINES_CONFIG_LANE_ARBITER_NUM_MEMORY   (ENGINES_CONFIG_LANE_ARBITER_NUM_MEMORY    ),
.ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST  (ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_REQUEST   ),
.ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE  (ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_CONTROL_RESPONSE ),
.ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE   (ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_ENGINE    ),
.ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY   (ENGINES_CONFIG_LANE_FIFO_ARBITER_SIZE_MEMORY    ),
.ENGINES_CONFIG_MAX_CAST_WIDTH_ARRAY     (ENGINES_CONFIG_MAX_CAST_WIDTH_ARRAY              ),
.ENGINES_CONFIG_MAX_MERGE_WIDTH_ARRAY    (ENGINES_CONFIG_MAX_MERGE_WIDTH_ARRAY             ),
.ENGINES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY (ENGINES_CONFIG_MERGE_CONNECT_PREFIX_ARRAY      ),
.ENGINES_COUNT_ARRAY                     (ENGINES_COUNT_ARRAY                              ),
.ENGINES_ENGINE_ID_ARRAY                 (ENGINES_ENGINE_ID_ARRAY                          ),
.ID_CU                                   (ID_CU                                            ),
.NUM_BUNDLES                             (NUM_BUNDLES_MAX                                  ),
.NUM_ENGINES                             (NUM_ENGINES                                      ),
.NUM_BACKTRACK_LANES                     (NUM_BACKTRACK_LANES                              ),
.NUM_LANES                               (NUM_LANES                                        )


