.ID_CU                               (ID_CU                               ),
.ID_BUNDLE                           (i                                   ),
.NUM_BUNDLES                         (NUM_BUNDLES                         ),
.NUM_LANES                           (LANES_COUNT_ARRAY[i]                ),
.NUM_ENGINES                         (NUM_ENGINES                         ),
.LANES_COUNT_ARRAY                   (LANES_COUNT_ARRAY                   ),
.ENGINES_COUNT_ARRAY                 (LANES_ENGINES_COUNT_ARRAY[i]        ),
.LANES_ENGINES_COUNT_ARRAY           (LANES_ENGINES_COUNT_ARRAY           ),
.ENGINES_CONFIG_ARRAY                (ENGINES_CONFIG_ARRAY                ),
.ENGINES_ENGINE_ID_ARRAY             (ENGINES_ENGINE_ID_ARRAY             ),
.LANES_CONFIG_ARRAY                  (BUNDLES_CONFIG_ARRAY[i]             ),
.BUNDLES_CONFIG_ARRAY                (BUNDLES_CONFIG_ARRAY                ),
.LANES_ENGINE_ID_ARRAY               (BUNDLES_ENGINE_ID_ARRAY[i]          ),
.BUNDLES_ENGINE_ID_ARRAY             (BUNDLES_ENGINE_ID_ARRAY             ),
.CU_BUNDLES_COUNT_ARRAY              (CU_BUNDLES_COUNT_ARRAY              ),
.CU_BUNDLES_LANES_COUNT_ARRAY        (CU_BUNDLES_LANES_COUNT_ARRAY        ),
.CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY(CU_BUNDLES_LANES_ENGINES_COUNT_ARRAY),
.CU_BUNDLES_CONFIG_ARRAY             (CU_BUNDLES_CONFIG_ARRAY             ),
.CU_BUNDLES_ENGINE_ID_ARRAY          (CU_BUNDLES_ENGINE_ID_ARRAY          ),

.LANES_CONFIG_MERGE_WIDTH_ARRAY      (BUNDLES_CONFIG_MERGE_WIDTH_ARRAY[i]          ),
.LANES_CONFIG_LANE_MERGE_WIDTH_ARRAY (BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY[i]     ),
.LANES_CONFIG_CAST_WIDTH_ARRAY       (BUNDLES_CONFIG_CAST_WIDTH_ARRAY[i]           ),
.LANES_CONFIG_LANE_CAST_WIDTH_ARRAY  (BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY[i]      ),
.LANES_CONFIG_MERGE_CONNECT_ARRAY    (BUNDLES_CONFIG_MERGE_CONNECT_ARRAY[i]        ),

.BUNDLES_CONFIG_MERGE_WIDTH_ARRAY      (BUNDLES_CONFIG_MERGE_WIDTH_ARRAY          ),
.BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY (BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY     ),
.BUNDLES_CONFIG_CAST_WIDTH_ARRAY       (BUNDLES_CONFIG_CAST_WIDTH_ARRAY           ),
.BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY  (BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY      ),
.BUNDLES_CONFIG_MERGE_CONNECT_ARRAY    (BUNDLES_CONFIG_MERGE_CONNECT_ARRAY        ),

.CU_BUNDLES_CONFIG_MERGE_WIDTH_ARRAY      (CU_BUNDLES_CONFIG_MERGE_WIDTH_ARRAY     ),
.CU_BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY (CU_BUNDLES_CONFIG_LANE_MERGE_WIDTH_ARRAY),
.CU_BUNDLES_CONFIG_CAST_WIDTH_ARRAY       (CU_BUNDLES_CONFIG_CAST_WIDTH_ARRAY      ),
.CU_BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY  (CU_BUNDLES_CONFIG_LANE_CAST_WIDTH_ARRAY ),
.CU_BUNDLES_CONFIG_MERGE_CONNECT_ARRAY    (CU_BUNDLES_CONFIG_MERGE_CONNECT_ARRAY   )