parameter NUM_CUS     = 1;
parameter NUM_BUNDLES = 4;
parameter NUM_LANES   = 4;
parameter NUM_ENGINES = 2;
parameter NUM_MODULES = 3;
parameter NUM_CUS_WIDTH_BITS     = 1;
parameter NUM_BUNDLES_WIDTH_BITS = 4;
parameter NUM_LANES_WIDTH_BITS   = 4;
parameter NUM_ENGINES_WIDTH_BITS = 2;
parameter NUM_MODULES_WIDTH_BITS = 3;
parameter CU_PACKET_SEQUENCE_ID_WIDTH_BITS = $clog2((192*NUM_BUNDLES)+(16*NUM_BUNDLES));
