
.m00_axi_read_in(kernel_s00_axi_read_out),
.m00_axi_read_out(kernel_s00_axi_read_in),
.m00_axi_write_in(kernel_s00_axi_write_out),
.m00_axi_write_out(kernel_s00_axi_write_in),
    

.m01_axi_read_in(kernel_s01_axi_read_out),
.m01_axi_read_out(kernel_s01_axi_read_in),
.m01_axi_write_in(kernel_s01_axi_write_out),
.m01_axi_write_out(kernel_s01_axi_write_in),
    