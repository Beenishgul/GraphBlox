parameter NUM_MEMORY_REQUESTOR = 2,
parameter ID_CU = 0,
// --------------------------------------------------------------------------------------
// CU SETTINGS
// --------------------------------------------------------------------------------------
`include "shared_parameters.vh"