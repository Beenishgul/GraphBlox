`include "global_timescale.vh"

import PKG_AXI4_FE::*;
import PKG_AXI4_MID::*;
import PKG_AXI4_BE::*;
import PKG_GLOBALS::*;
import PKG_CACHE::*;
import PKG_CONTROL::*;
import PKG_DESCRIPTOR::*;
import PKG_FUNCTIONS::*;
import PKG_MEMORY::*;
import PKG_ENGINE::*;
import PKG_SETUP::*;

