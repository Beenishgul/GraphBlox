    parameter ID_CU     = 0,
    parameter ID_BUNDLE = 0,
    parameter ID_LANE   = 0,
// --------------------------------------------------------------------------------------
// CU SETTINGS
// --------------------------------------------------------------------------------------
`include "shared_parameters.vh"

