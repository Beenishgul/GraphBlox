// -----------------------------------------------------------------------------
//
//    "GLay: A Vertex Centric Re-Configurable Graph Processing Overlay"
//
// -----------------------------------------------------------------------------
// Copyright (c) 2021-2023 All rights reserved
// -----------------------------------------------------------------------------
// Author : Abdullah Mughrabi atmughrabi@gmail.com/atmughra@virginia.edu
// File   : kernel_afu.sv
// Create : 2022-11-29 12:42:56
// Revise : 2023-06-13 00:31:13
// Editor : sublime text4, tab size (2)
// -----------------------------------------------------------------------------

`include "global_package.vh"

module kernel_afu (
  // System Signals
  input  logic                         ap_clk         ,
  input  logic                         ap_rst_n       ,
  // AXI4 master interface m00_axi
  output logic                         m00_axi_awvalid,
  input  logic                         m00_axi_awready,
  output logic [ M_AXI4_BE_ADDR_W-1:0] m00_axi_awaddr ,
  output logic [  M_AXI4_BE_LEN_W-1:0] m00_axi_awlen  ,
  output logic                         m00_axi_wvalid ,
  input  logic                         m00_axi_wready ,
  output logic [ M_AXI4_BE_DATA_W-1:0] m00_axi_wdata  ,
  output logic [ M_AXI4_BE_STRB_W-1:0] m00_axi_wstrb  ,
  output logic                         m00_axi_wlast  ,
  input  logic                         m00_axi_bvalid ,
  output logic                         m00_axi_bready ,
  output logic                         m00_axi_arvalid,
  input  logic                         m00_axi_arready,
  output logic [ M_AXI4_BE_ADDR_W-1:0] m00_axi_araddr ,
  output logic [  M_AXI4_BE_LEN_W-1:0] m00_axi_arlen  ,
  input  logic                         m00_axi_rvalid ,
  output logic                         m00_axi_rready ,
  input  logic [ M_AXI4_BE_DATA_W-1:0] m00_axi_rdata  ,
  input  logic                         m00_axi_rlast  ,
  // Control Signals
  // AXI4 master interface m00_axi missing ports
  input  logic [   M_AXI4_BE_ID_W-1:0] m00_axi_bid    ,
  input  logic [   M_AXI4_BE_ID_W-1:0] m00_axi_rid    ,
  input  logic [ M_AXI4_BE_RESP_W-1:0] m00_axi_rresp  ,
  input  logic [ M_AXI4_BE_RESP_W-1:0] m00_axi_bresp  ,
  output logic [   M_AXI4_BE_ID_W-1:0] m00_axi_awid   ,
  output logic [ M_AXI4_BE_SIZE_W-1:0] m00_axi_awsize ,
  output logic [M_AXI4_BE_BURST_W-1:0] m00_axi_awburst,
  output logic [ M_AXI4_BE_LOCK_W-1:0] m00_axi_awlock ,
  output logic [M_AXI4_BE_CACHE_W-1:0] m00_axi_awcache,
  output logic [ M_AXI4_BE_PROT_W-1:0] m00_axi_awprot ,
  output logic [  M_AXI4_BE_QOS_W-1:0] m00_axi_awqos  ,
  output logic [   M_AXI4_BE_ID_W-1:0] m00_axi_arid   ,
  output logic [ M_AXI4_BE_SIZE_W-1:0] m00_axi_arsize ,
  output logic [M_AXI4_BE_BURST_W-1:0] m00_axi_arburst,
  output logic [ M_AXI4_BE_LOCK_W-1:0] m00_axi_arlock ,
  output logic [M_AXI4_BE_CACHE_W-1:0] m00_axi_arcache,
  output logic [ M_AXI4_BE_PROT_W-1:0] m00_axi_arprot ,
  output logic [  M_AXI4_BE_QOS_W-1:0] m00_axi_arqos  ,
  input  logic                         ap_start       ,
  output logic                         ap_idle        ,
  output logic                         ap_done        ,
  output logic                         ap_ready       ,
  input  logic                         ap_continue    ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_0       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_1       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_2       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_3       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_4       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_5       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_6       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_7       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_8       ,
  input  logic [ M_AXI4_BE_ADDR_W-1:0] buffer_9
);

genvar i;
// --------------------------------------------------------------------------------------
// Wires and Variables
// --------------------------------------------------------------------------------------
logic areset_m_axi  ;
logic areset_cu     ;
logic areset_control;


logic endian_read_reg ;
logic endian_write_reg;

// --------------------------------------------------------------------------------------
// Kernel -> State Control
// --------------------------------------------------------------------------------------
ControlChainInterfaceInput  kernel_control_in ;
ControlChainInterfaceOutput kernel_control_out;

KernelDescriptorPayload kernel_control_descriptor_in ;
KernelDescriptor        kernel_control_descriptor_out;

logic kernel_cu_done_out         ;
logic kernel_cu_fifo_setup_signal;

// --------------------------------------------------------------------------------------
// CU -> [CU_CACHE|BUNDLES|LANES|ENGINES]
// --------------------------------------------------------------------------------------
KernelDescriptor kernel_cu_descriptor_in;

// --------------------------------------------------------------------------------------
// System Cache -> AXI Mutli channels support
// --------------------------------------------------------------------------------------
logic areset_axi_slice[GLOBAL_NUM_CHANNELS-1:0];
logic areset_cache    [GLOBAL_NUM_CHANNELS-1:0];
// --------------------------------------------------------------------------------------
// AXI
// --------------------------------------------------------------------------------------
AXI4BEMasterReadInterface  m_axi4_read [GLOBAL_NUM_CHANNELS-1:0];
AXI4BEMasterWriteInterface m_axi4_write[GLOBAL_NUM_CHANNELS-1:0];

AXI4MIDSlaveReadInterfaceOutput  kernel_s_axi_read_out [GLOBAL_NUM_CHANNELS-1:0];
AXI4MIDSlaveReadInterfaceInput   kernel_s_axi_read_in  [GLOBAL_NUM_CHANNELS-1:0];
AXI4MIDSlaveWriteInterfaceOutput kernel_s_axi_write_out[GLOBAL_NUM_CHANNELS-1:0];
AXI4MIDSlaveWriteInterfaceInput  kernel_s_axi_write_in [GLOBAL_NUM_CHANNELS-1:0];

AXI4BEMasterReadInterfaceInput   kernel_m_axi4_read_in  [GLOBAL_NUM_CHANNELS-1:0];
AXI4BEMasterReadInterfaceOutput  kernel_m_axi4_read_out [GLOBAL_NUM_CHANNELS-1:0];
AXI4BEMasterWriteInterfaceInput  kernel_m_axi4_write_in [GLOBAL_NUM_CHANNELS-1:0];
AXI4BEMasterWriteInterfaceOutput kernel_m_axi4_write_out[GLOBAL_NUM_CHANNELS-1:0];

logic [GLOBAL_NUM_CHANNELS-1:0] kernel_cache_setup_signal;

// --------------------------------------------------------------------------------------
//   Register and invert reset signal.
// --------------------------------------------------------------------------------------
parameter PULSE_HOLD    = 100;
logic     areset_system      ;
// --------------------------------------------------------------------------------------
always_ff @(posedge ap_clk) begin
  areset_m_axi   <= areset_system;
  areset_cu      <= areset_system;
  areset_control <= areset_system;

  for (int i = 0; i < GLOBAL_NUM_CHANNELS; i++) begin
    areset_cache[i]     <= areset_system;
    areset_axi_slice[i] <= areset_system;
  end
end

logic [PULSE_HOLD-1:0] sync_ff;

always_ff @(posedge ap_clk or negedge ap_rst_n) begin
  if (~ap_rst_n | ap_done) begin
    // Asynchronously assert reset (active low reset)
    sync_ff <= {PULSE_HOLD{1'b1}};;
  end else begin
    // Synchronously de-assert reset
    sync_ff <= sync_ff << 1'b1;
  end
end

// Output of the second flip-flop is the synchronized reset
assign areset_system = sync_ff[PULSE_HOLD-1];

// --------------------------------------------------------------------------------------
// Control chain signals
// --------------------------------------------------------------------------------------
always_ff @(posedge ap_clk) begin
  if (areset_control) begin
    kernel_control_in.ap_start    <= 1'b0;
    kernel_control_in.ap_continue <= 1'b0;
    kernel_control_in.setup       <= 1'b0;
    kernel_control_in.done        <= 1'b0;
  end
  else begin
    kernel_control_in.ap_start    <= ap_start;
    kernel_control_in.ap_continue <= ap_continue;
    kernel_control_in.setup       <= ~(kernel_cu_fifo_setup_signal | (|kernel_cache_setup_signal));
    kernel_control_in.done        <= kernel_cu_done_out;
  end
end

always_ff @(posedge ap_clk) begin
  if (areset_control) begin
    ap_ready         <= 1'b0;
    ap_done          <= 1'b0;
    ap_idle          <= 1'b1;
    endian_read_reg  <= 1'b0;
    endian_write_reg <= 1'b0;
  end
  else begin
    ap_done          <= kernel_control_out.ap_done;
    ap_ready         <= kernel_control_out.ap_ready;
    ap_idle          <= kernel_control_out.ap_idle;
    endian_read_reg  <= kernel_control_out.endian_read;
    endian_write_reg <= kernel_control_out.endian_write;
  end
end

// --------------------------------------------------------------------------------------
// READ AXI4 SIGNALS INPUT
// --------------------------------------------------------------------------------------
assign m_axi4_read[0].in.rvalid  = m00_axi_rvalid ; // Read channel valid
assign m_axi4_read[0].in.arready = m00_axi_arready; // Address read channel ready
assign m_axi4_read[0].in.rlast   = m00_axi_rlast  ; // Read channel last word
assign m_axi4_read[0].in.rdata   = swap_endianness_cacheline_axi_be(m00_axi_rdata, endian_read_reg)  ; // Read channel data
assign m_axi4_read[0].in.rid     = m00_axi_rid    ; // Read channel ID
assign m_axi4_read[0].in.rresp   = m00_axi_rresp  ; // Read channel response


// --------------------------------------------------------------------------------------
// READ AXI4 SIGNALS OUTPUT
// --------------------------------------------------------------------------------------
assign m00_axi_arvalid = m_axi4_read[0].out.arvalid; // Address read channel valid
assign m00_axi_araddr  = m_axi4_read[0].out.araddr ; // Address read channel address
assign m00_axi_arlen   = m_axi4_read[0].out.arlen  ; // Address write channel burst length
assign m00_axi_rready  = m_axi4_read[0].out.rready ; // Read channel ready
assign m00_axi_arid    = m_axi4_read[0].out.arid   ; // Address read channel ID
assign m00_axi_arsize  = m_axi4_read[0].out.arsize ; // Address read channel burst size. This signal indicates the size of each transfer in the burst
assign m00_axi_arburst = m_axi4_read[0].out.arburst; // Address read channel burst type
assign m00_axi_arlock  = m_axi4_read[0].out.arlock ; // Address read channel lock type
assign m00_axi_arcache = m_axi4_read[0].out.arcache; // Address read channel memory type. Transactions set with Normal Non-cacheable Modifiable and Bufferable (0011).
assign m00_axi_arprot  = m_axi4_read[0].out.arprot ; // Address write channel protection type. Transactions set with Normal, Secure, and Data attributes (000).
assign m00_axi_arqos   = m_axi4_read[0].out.arqos  ; // Address write channel quality of service


// --------------------------------------------------------------------------------------
// WRITE AXI4 SIGNALS INPUT
// --------------------------------------------------------------------------------------
assign m_axi4_write[0].in.awready = m00_axi_awready; // Address write channel ready
assign m_axi4_write[0].in.wready  = m00_axi_wready ; // Write channel ready
assign m_axi4_write[0].in.bid     = m00_axi_bid    ; // Write response channel ID
assign m_axi4_write[0].in.bresp   = m00_axi_bresp  ; // Write channel response
assign m_axi4_write[0].in.bvalid  = m00_axi_bvalid ; // Write response channel valid


// --------------------------------------------------------------------------------------
// WRITE AXI4 SIGNALS OUTPUT
// --------------------------------------------------------------------------------------
assign m00_axi_awvalid = m_axi4_write[0].out.awvalid; // Address write channel valid
assign m00_axi_awid    = m_axi4_write[0].out.awid   ; // Address write channel ID
assign m00_axi_awaddr  = m_axi4_write[0].out.awaddr ; // Address write channel address
assign m00_axi_awlen   = m_axi4_write[0].out.awlen  ; // Address write channel burst length
assign m00_axi_awsize  = m_axi4_write[0].out.awsize ; // Address write channel burst size. This signal indicates the size of each transfer in the burst
assign m00_axi_awburst = m_axi4_write[0].out.awburst; // Address write channel burst type
assign m00_axi_awlock  = m_axi4_write[0].out.awlock ; // Address write channel lock type
assign m00_axi_awcache = m_axi4_write[0].out.awcache; // Address write channel memory type. Transactions set with Normal Non-cacheable Modifiable and Bufferable (0011).
assign m00_axi_awprot  = m_axi4_write[0].out.awprot ; // Address write channel protection type. Transactions set with Normal, Secure, and Data attributes (000).
assign m00_axi_awqos   = m_axi4_write[0].out.awqos  ; // Address write channel quality of service
assign m00_axi_wdata   = swap_endianness_cacheline_axi_be(m_axi4_write[0].out.wdata , endian_write_reg); // Write channel data
assign m00_axi_wstrb   = m_axi4_write[0].out.wstrb  ; // Write channel write strobe
assign m00_axi_wlast   = m_axi4_write[0].out.wlast  ; // Write channel last word flag
assign m00_axi_wvalid  = m_axi4_write[0].out.wvalid ; // Write channel valid
assign m00_axi_bready  = m_axi4_write[0].out.bready ; // Write response channel ready

// --------------------------------------------------------------------------------------
// DRIVE DESCRIPTOR
// --------------------------------------------------------------------------------------
always_ff @(posedge ap_clk) begin
  kernel_control_descriptor_in.buffer_0 <= buffer_0  ;
  kernel_control_descriptor_in.buffer_1 <= buffer_1  ;
  kernel_control_descriptor_in.buffer_2 <= buffer_2  ;
  kernel_control_descriptor_in.buffer_3 <= buffer_3  ;
  kernel_control_descriptor_in.buffer_4 <= buffer_4  ;
  kernel_control_descriptor_in.buffer_5 <= buffer_5  ;
  kernel_control_descriptor_in.buffer_6 <= buffer_6  ;
  kernel_control_descriptor_in.buffer_7 <= buffer_7  ;
  kernel_control_descriptor_in.buffer_8 <= buffer_8  ;
  kernel_control_descriptor_in.buffer_9 <= buffer_9  ;
end


generate
  if(GLOBAL_SYSTEM_CACHE_IP == 1) begin
// --------------------------------------------------------------------------------------
// System Cache CH 0-> AXI
// --------------------------------------------------------------------------------------
    kernel_cache inst_kernel_cache_ch0 (
      .ap_clk            (ap_clk                      ),
      .areset            (areset_cache[0]             ),
      .s_axi_read_out    (kernel_s_axi_read_out[0]    ),
      .s_axi_read_in     (kernel_s_axi_read_in[0]     ),
      .s_axi_write_out   (kernel_s_axi_write_out[0]   ),
      .s_axi_write_in    (kernel_s_axi_write_in[0]    ),
      .m_axi_read_in     (kernel_m_axi4_read_in[0]    ),
      .m_axi_read_out    (kernel_m_axi4_read_out[0]   ),
      .m_axi_write_in    (kernel_m_axi4_write_in[0]   ),
      .m_axi_write_out   (kernel_m_axi4_write_out[0]  ),
      .cache_setup_signal(kernel_cache_setup_signal[0])
    );
  end else begin
    assign kernel_cache_setup_signal[0] = 0;
    assign kernel_s_axi_read_out[0]     = kernel_m_axi4_read_in[0];
    assign kernel_m_axi4_read_out[0]    = kernel_s_axi_read_in[0];
    assign kernel_s_axi_write_out[0]    = kernel_m_axi4_write_in[0];
    assign kernel_m_axi4_write_out[0]   = kernel_s_axi_write_in[0];
  end
endgenerate

generate
  if(GLOBAL_NUM_CHANNELS > 1) begin
    if(GLOBAL_SYSTEM_STREAM_IP == 1) begin
// --------------------------------------------------------------------------------------
// System Cache CH 1 -> AXI
// --------------------------------------------------------------------------------------
      kernel_cache inst_kernel_cache_ch1 (
        .ap_clk            (ap_clk                      ),
        .areset            (areset_cache[1]             ),
        .s_axi_read_out    (kernel_s_axi_read_out[1]    ),
        .s_axi_read_in     (kernel_s_axi_read_in[1]     ),
        .s_axi_write_out   (kernel_s_axi_write_out[1]   ),
        .s_axi_write_in    (kernel_s_axi_write_in[1]    ),
        .m_axi_read_in     (kernel_m_axi4_read_in[1]    ),
        .m_axi_read_out    (kernel_m_axi4_read_out[1]   ),
        .m_axi_write_in    (kernel_m_axi4_write_in[1]   ),
        .m_axi_write_out   (kernel_m_axi4_write_out[1]  ),
        .cache_setup_signal(kernel_cache_setup_signal[1])
      );
    end else begin
      assign kernel_cache_setup_signal[1] = 0;
      assign kernel_s_axi_read_out[1]     = kernel_m_axi4_read_in[1];
      assign kernel_m_axi4_read_out[1]    = kernel_s_axi_read_in[1];
      assign kernel_s_axi_write_out[1]    = kernel_m_axi4_write_in[1];
      assign kernel_m_axi4_write_out[1]   = kernel_s_axi_write_in[1];
    end
  end
endgenerate

// --------------------------------------------------------------------------------------
// Kernel CACHE (M->S) Register Slice
// --------------------------------------------------------------------------------------
// --------------------------------------------------------------------------------------
generate
  for (i=0; i<(GLOBAL_NUM_CHANNELS); i++) begin : generate_axi_register_slice_be_ch
// --------------------------------------------------------------------------------------
    axi_register_slice_back_end inst_axi_register_slice_be (
      .ap_clk         (ap_clk                    ),
      .areset         (areset_axi_slice[i]       ),
      .s_axi_read_out (kernel_m_axi4_read_in[i]  ),
      .s_axi_read_in  (kernel_m_axi4_read_out[i] ),
      .s_axi_write_out(kernel_m_axi4_write_in[i] ),
      .s_axi_write_in (kernel_m_axi4_write_out[i]),
      .m_axi_read_in  (m_axi4_read[i].in         ),
      .m_axi_read_out (m_axi4_read[i].out        ),
      .m_axi_write_in (m_axi4_write[i].in        ),
      .m_axi_write_out(m_axi4_write[i].out       )
    );
  end
endgenerate

// --------------------------------------------------------------------------------------
// CU -> [CU_CACHE|BUNDLES|LANES|ENGINES]
// --------------------------------------------------------------------------------------
// Kernel_setup
assign kernel_cu_descriptor_in = kernel_control_descriptor_out;

kernel_cu #(
  .ID_CU       (0                  ),
  .NUM_CHANNELS(GLOBAL_NUM_CHANNELS)
) inst_kernel_cu (
  .ap_clk           (ap_clk                     ),
  .areset           (areset_cu                  ),
  .descriptor_in    (kernel_cu_descriptor_in    ),
  .m_axi_read_in    (kernel_s_axi_read_out      ),
  .m_axi_read_out   (kernel_s_axi_read_in       ),
  .m_axi_write_in   (kernel_s_axi_write_out     ),
  .m_axi_write_out  (kernel_s_axi_write_in      ),
  .fifo_setup_signal(kernel_cu_fifo_setup_signal),
  .done_out         (kernel_cu_done_out         )
);

// --------------------------------------------------------------------------------------
// Kernel -> State Control
// --------------------------------------------------------------------------------------
kernel_control inst_kernel_control (
  .ap_clk        (ap_clk                       ),
  .areset        (areset_control               ),
  .control_in    (kernel_control_in            ),
  .control_out   (kernel_control_out           ),
  .descriptor_in (kernel_control_descriptor_in ),
  .descriptor_out(kernel_control_descriptor_out)
);

endmodule : kernel_afu

