
        .C_M00_AXI_ADDR_WIDTH      (C_M00_AXI_ADDR_WIDTH      ),
        .C_M00_AXI_DATA_WIDTH      (C_M00_AXI_DATA_WIDTH      ),
        

        .C_M01_AXI_ADDR_WIDTH      (C_M01_AXI_ADDR_WIDTH      ),
        .C_M01_AXI_DATA_WIDTH      (C_M01_AXI_DATA_WIDTH      ),
        